//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9 (64-bit)
//Part Number: GW5A-LV25MG121NES
//Device: GW5A-25
//Device Version: A
//Created Time: Sat Apr 20 11:36:50 2024

module blk_mem_gen_0 (dout, clk, oce, ce, reset, wre, ad, din, byte_en);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [13:0] ad;
input [31:0] din;
input [3:0] byte_en;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire [15:0] sp_inst_0_dout_w;
wire [15:0] sp_inst_0_dout;
wire [15:0] sp_inst_1_dout_w;
wire [15:0] sp_inst_1_dout;
wire [15:0] sp_inst_2_dout_w;
wire [15:0] sp_inst_2_dout;
wire [15:0] sp_inst_3_dout_w;
wire [15:0] sp_inst_3_dout;
wire [15:0] sp_inst_4_dout_w;
wire [15:0] sp_inst_4_dout;
wire [15:0] sp_inst_5_dout_w;
wire [15:0] sp_inst_5_dout;
wire [15:0] sp_inst_6_dout_w;
wire [15:0] sp_inst_6_dout;
wire [15:0] sp_inst_7_dout_w;
wire [15:0] sp_inst_7_dout;
wire [15:0] sp_inst_8_dout_w;
wire [15:0] sp_inst_8_dout;
wire [15:0] sp_inst_9_dout_w;
wire [15:0] sp_inst_9_dout;
wire [15:0] sp_inst_10_dout_w;
wire [15:0] sp_inst_10_dout;
wire [15:0] sp_inst_11_dout_w;
wire [15:0] sp_inst_11_dout;
wire [15:0] sp_inst_12_dout_w;
wire [15:0] sp_inst_12_dout;
wire [15:0] sp_inst_13_dout_w;
wire [15:0] sp_inst_13_dout;
wire [15:0] sp_inst_14_dout_w;
wire [15:0] sp_inst_14_dout;
wire [15:0] sp_inst_15_dout_w;
wire [15:0] sp_inst_15_dout;
wire [15:0] sp_inst_16_dout_w;
wire [31:16] sp_inst_16_dout;
wire [15:0] sp_inst_17_dout_w;
wire [31:16] sp_inst_17_dout;
wire [15:0] sp_inst_18_dout_w;
wire [31:16] sp_inst_18_dout;
wire [15:0] sp_inst_19_dout_w;
wire [31:16] sp_inst_19_dout;
wire [15:0] sp_inst_20_dout_w;
wire [31:16] sp_inst_20_dout;
wire [15:0] sp_inst_21_dout_w;
wire [31:16] sp_inst_21_dout;
wire [15:0] sp_inst_22_dout_w;
wire [31:16] sp_inst_22_dout;
wire [15:0] sp_inst_23_dout_w;
wire [31:16] sp_inst_23_dout;
wire [15:0] sp_inst_24_dout_w;
wire [31:16] sp_inst_24_dout;
wire [15:0] sp_inst_25_dout_w;
wire [31:16] sp_inst_25_dout;
wire [15:0] sp_inst_26_dout_w;
wire [31:16] sp_inst_26_dout;
wire [15:0] sp_inst_27_dout_w;
wire [31:16] sp_inst_27_dout;
wire [15:0] sp_inst_28_dout_w;
wire [31:16] sp_inst_28_dout;
wire [15:0] sp_inst_29_dout_w;
wire [31:16] sp_inst_29_dout;
wire [15:0] sp_inst_30_dout_w;
wire [31:16] sp_inst_30_dout;
wire [15:0] sp_inst_31_dout_w;
wire [31:16] sp_inst_31_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_60;
wire mux_o_61;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_123;
wire mux_o_124;
wire mux_o_125;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_154;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_245;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_251;
wire mux_o_252;
wire mux_o_253;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_258;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_265;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_270;
wire mux_o_271;
wire mux_o_272;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_278;
wire mux_o_279;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_308;
wire mux_o_309;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_321;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_335;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_349;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_356;
wire mux_o_357;
wire mux_o_358;
wire mux_o_360;
wire mux_o_361;
wire mux_o_362;
wire mux_o_363;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_370;
wire mux_o_371;
wire mux_o_372;
wire mux_o_373;
wire mux_o_375;
wire mux_o_376;
wire mux_o_377;
wire mux_o_378;
wire mux_o_379;
wire mux_o_380;
wire mux_o_381;
wire mux_o_382;
wire mux_o_383;
wire mux_o_384;
wire mux_o_385;
wire mux_o_386;
wire mux_o_387;
wire mux_o_388;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_401;
wire mux_o_402;
wire mux_o_403;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_408;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_412;
wire mux_o_413;
wire mux_o_414;
wire mux_o_415;
wire mux_o_416;
wire mux_o_417;
wire mux_o_418;
wire mux_o_420;
wire mux_o_421;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_426;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_431;
wire mux_o_432;
wire mux_o_433;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_440;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_453;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_460;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_465;
wire mux_o_466;
wire mux_o_467;
wire mux_o_468;
wire mux_o_469;
wire mux_o_470;
wire mux_o_471;
wire mux_o_472;
wire mux_o_473;
wire mux_o_474;
wire mux_o_475;
wire mux_o_476;
wire mux_o_477;
wire mux_o_478;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_0.INIT = 16'h0001;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_1.INIT = 16'h0002;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_2.INIT = 16'h0004;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_3.INIT = 16'h0008;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_4.INIT = 16'h0010;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_5.INIT = 16'h0020;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_6.INIT = 16'h0040;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_7.INIT = 16'h0080;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_8.INIT = 16'h0100;
LUT4 lut_inst_9 (
  .F(lut_f_9),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_9.INIT = 16'h0200;
LUT4 lut_inst_10 (
  .F(lut_f_10),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_10.INIT = 16'h0400;
LUT4 lut_inst_11 (
  .F(lut_f_11),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_11.INIT = 16'h0800;
LUT4 lut_inst_12 (
  .F(lut_f_12),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_12.INIT = 16'h1000;
LUT4 lut_inst_13 (
  .F(lut_f_13),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_13.INIT = 16'h2000;
LUT4 lut_inst_14 (
  .F(lut_f_14),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_14.INIT = 16'h4000;
LUT4 lut_inst_15 (
  .F(lut_f_15),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_15.INIT = 16'h8000;
SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[15:0],sp_inst_0_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b01;
defparam sp_inst_0.BIT_WIDTH = 16;
defparam sp_inst_0.BLK_SEL = 3'b001;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h000CD1CF358E31EF002F018C002C11AD020F3590020F35F0B1EF012F2000000D;
defparam sp_inst_0.INIT_RAM_01 = 256'hFD8CE3EC118CFD8C002C102C000C302C002CF9AC118C018011AC01AD000D018C;
defparam sp_inst_0.INIT_RAM_02 = 256'h0000000000000000002080000020B000F06300230180200C402C418CA06C442C;
defparam sp_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[15:0],sp_inst_1_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_1}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b01;
defparam sp_inst_1.BIT_WIDTH = 16;
defparam sp_inst_1.BLK_SEL = 3'b001;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'h92A8A2A7B2A6C2A5D2A472B482B392B2A2B1B2B0C2AFD2AEE2ADF2AC0055C435;
defparam sp_inst_1.INIT_RAM_01 = 256'h2DA0818D2DA0418D2DA0218D2DA0118D65A0F18D140C42A352A162AB72AA82A9;
defparam sp_inst_1.INIT_RAM_02 = 256'h1400B8001C00B000240098002C0064003400E0003C00A0002DA0018D2DA0018D;
defparam sp_inst_1.INIT_RAM_03 = 256'hC2A5D2A472B482B392B2A2B1B2B0C2AFD2AEE2ADF2AC0055040050000DA0018D;
defparam sp_inst_1.INIT_RAM_04 = 256'h0184D00CF51F81081508D0083800C41542A352A162AB72AA82A992A8A2A7B2A6;
defparam sp_inst_1.INIT_RAM_05 = 256'hAFFF02040190198CBD8CB4AC2DC00085700F200E000DE0C600060061F0630020;
defparam sp_inst_1.INIT_RAM_06 = 256'hF51F81081508D0082580012C008900201063006197FF2804DBFFFDCEF1EF91AD;
defparam sp_inst_1.INIT_RAM_07 = 256'hB2B0C2AFD2AEE2ADF2AC0055C4350020F51F01081508D008DFFF052900ECD007;
defparam sp_inst_1.INIT_RAM_08 = 256'hB2A6C2A5D2A4E2BFF2BE02BD12BC22BB32BA42B952B862B772B482B392B2A2B1;
defparam sp_inst_1.INIT_RAM_09 = 256'h058CF1ACD60D00001195C41502AC22B632A242A352A162AB72AA82A992A8A2A7;
defparam sp_inst_1.INIT_RAM_0A = 256'h72B482B392B2A2B1B2B0C2AFD2AEE2ADF2AC005513FFF08400048000F1ACF99F;
defparam sp_inst_1.INIT_RAM_0B = 256'h72AA82A992A8A2A7B2A6C2A5D2A4E2BFF2BE02BD12BC22BB32BA42B952B862B7;
defparam sp_inst_1.INIT_RAM_0C = 256'h00AC72C4C076B07640630020C40C018C100CC42C12B522B632A242A352A162AB;
defparam sp_inst_1.INIT_RAM_0D = 256'hAECC4D80058C31ACAECC6ACD6C00AEC0B2CC018C72CC82C0B2C092C06ACC52C6;
defparam sp_inst_1.INIT_RAM_0E = 256'h31ACB2CD31AC92CC52CDB2CCB1ACB2CD300C82CC82CC31AC92CC0C0D92CC858C;
defparam sp_inst_1.INIT_RAM_0F = 256'hB07640630020C063B0760000018DB2CD72CC918D3C0CAECDAECC058CAECCB2CC;
defparam sp_inst_1.INIT_RAM_10 = 256'hB2CD62CCB2CC058CB2CC098D01ADCE0C31ADB2CC72CD2800B2C062C572C4C076;
defparam sp_inst_1.INIT_RAM_11 = 256'h018D81AD09AD31CCB2CC72CECE0D2C00B2C0F19F118C818C058CCE0C0000D5AC;
defparam sp_inst_1.INIT_RAM_12 = 256'h62CCCE0DF19F058C818C058CCE0C0000C98DB2CC018DFD8C62CCB2CC058CB2CC;
defparam sp_inst_1.INIT_RAM_13 = 256'hB2C062C572C4C076B07640630020C063B0760000018D81AD09AD31CC72CEFD8C;
defparam sp_inst_1.INIT_RAM_14 = 256'h00006800A2C0D58D0C0CB2CDB2CC058CB2CC098D01ADCE0C31ADB2CC72CD2800;
defparam sp_inst_1.INIT_RAM_15 = 256'hCE0C31ADB2CC72CD018D81AD09AD31CCA2CC72CECE0DF19F058C818C058CCE0C;
defparam sp_inst_1.INIT_RAM_16 = 256'h818C058CCE0C0000440095ACB2CD62CCA2CC058CA2CCB2CC058CB2CC098D01AD;
defparam sp_inst_1.INIT_RAM_17 = 256'h0000B9ACA2CD62CCA2CC058CA2CC018D81AD09AD31CCA2CC72CECE0DF19F058C;
defparam sp_inst_1.INIT_RAM_18 = 256'h818E158CCE0C158D81AD05ADCE0C818D158CCE0C40763076C0630020C063B076;
defparam sp_inst_1.INIT_RAM_19 = 256'hCE0C818D158CCE0C40763076C0630020406330760000158D81ADB5CDBC0DCE0C;
defparam sp_inst_1.INIT_RAM_1A = 256'h706180630020406330760000158D81AD41ADCE0C818D158CCE0C158D81AD05AD;
defparam sp_inst_1.INIT_RAM_1B = 256'h8063607670610184B6CC7FFF17FF01840805B2CC3BFFB2CC140CB2C080766076;
defparam sp_inst_1.INIT_RAM_1C = 256'h806300204063207630610000F59F058C008CA3FF0000407620763061C0630020;
defparam sp_inst_1.INIT_RAM_1D = 256'h607670610000F7FF8FFF01840405B2CCB3FFAFFFB2CC180CB2C0807660767061;
defparam sp_inst_1.INIT_RAM_1E = 256'h3FFF01841005B2CC63FFBEC0BAC0B6C0B2CC400C807660767061806300208063;
defparam sp_inst_1.INIT_RAM_1F = 256'hC076A076B061406300208063607670610184018CB2CC97FF2FFF01840805B2CC;
defparam sp_inst_1.INIT_RAM_20 = 256'h72CCA18C72CCBACC818C72CC72CCA18C72CCBECC818C72CCB2CC600CB2C072C4;
defparam sp_inst_1.INIT_RAM_21 = 256'h0020C063A076B06100009FFF03FF9BFF01841005B2CCBFFFF3FFB6CC818C72CC;
defparam sp_inst_1.INIT_RAM_22 = 256'h72CCA18C72CCBECC818C72CCB2CC080CB2C052C662C572C4C076A076B0614063;
defparam sp_inst_1.INIT_RAM_23 = 256'h52C503FF01841005B2CC27FF5BFFB6CC818C72CC72CCA18C72CCBACC818C72CC;
defparam sp_inst_1.INIT_RAM_24 = 256'h52C662C572C4C076A076B06140630020C063A076B0610000FBFF5FFFE7FF62C4;
defparam sp_inst_1.INIT_RAM_25 = 256'h72CC72CCA18C72CCBACC818C72CC72CCA18C72CCBECC818C72CCB2CC0C0CB2C0;
defparam sp_inst_1.INIT_RAM_26 = 256'h0020C063A076B0610000BFFF47FF62C452C563FF01841005B2CC87FFB6CC818C;
defparam sp_inst_1.INIT_RAM_27 = 256'h4063002080636076706100003C00D0040185BECCBECC008C8076607670618063;
defparam sp_inst_1.INIT_RAM_28 = 256'h87FFB40492CC300C72CC1D8072CC258042CC42C752C662C572C4C076A076B061;
defparam sp_inst_1.INIT_RAM_29 = 256'h52CDC1AC35CDC2CEB2CD5DCC00070980B1AE92CD52CC5000B2C092CC72CC0C00;
defparam sp_inst_1.INIT_RAM_2A = 256'h358CB5CE31ADB2CEB2CD62CCB19F92CCB2CC058CB2CC92CC000709A035CC92CE;
defparam sp_inst_1.INIT_RAM_2B = 256'h240C82CD82CC000C0800C18C31ACC2CDFD8CA2CC1D8DB2CCA2CD7400A2CC31CC;
defparam sp_inst_1.INIT_RAM_2C = 256'hA2CCA2CCFD8CA2CC97FF0184818C5D8C818C82CC1400818CC18C818C82CC198D;
defparam sp_inst_1.INIT_RAM_2D = 256'h0DAC280CBECD300072C4C076A076B06140630020C063A076B0610184000C8C0C;
defparam sp_inst_1.INIT_RAM_2E = 256'hB0610184000CC59FBECCBECC018C72CC72CC058C72CC33FF0184BECC3FFF3404;
defparam sp_inst_1.INIT_RAM_2F = 256'h82CC72CB62CA52C942C832C722C612C532C40076E076F06180630020C063A076;
defparam sp_inst_1.INIT_RAM_30 = 256'h92CC040CE5AC940C8ECD8ECC018C31AC32CDB2CC3000B2C0A2CC72CC72CC918C;
defparam sp_inst_1.INIT_RAM_31 = 256'h018CA2CC0180018C31ACE18C00CC898DADAC4C0D6D8C018C31AC32CD058CB2CC;
defparam sp_inst_1.INIT_RAM_32 = 256'h118CA2CC0FFF0184818C018CA2CC9800B2CC058CB2CCA2CC118CA2CCDBFF0184;
defparam sp_inst_1.INIT_RAM_33 = 256'hB2CCA2CC118CA2CC13FF018492C528060007018CA2CC6800B2CC058CB2CCA2CC;
defparam sp_inst_1.INIT_RAM_34 = 256'hB2CC058CB2CCA2CC118CA2CCDBFF018492C528060407018CA2CC3000B2CC058C;
defparam sp_inst_1.INIT_RAM_35 = 256'hA2CCC000B2CC058CB2CCA2CC118CA2CCA3FF018492C520060007018CA2CCF800;
defparam sp_inst_1.INIT_RAM_36 = 256'h0007018CA2CC8800B2CC058CB2CCA2CC118CA2CC6BFF018492C508060007018C;
defparam sp_inst_1.INIT_RAM_37 = 256'hB2CC058CB2CCD3FF94045000B2CC058CB2CCA2CC118CA2CC33FF018492C54006;
defparam sp_inst_1.INIT_RAM_38 = 256'h31AC418C018C31CC32CE058CB2CC31AD280C92CD3C0092C0B2CC058CB2CC3800;
defparam sp_inst_1.INIT_RAM_39 = 256'h018D31AC32CD058CB2CCD98DC00C018D31AC32CD058CB2CCB2CC058CB2CC92CC;
defparam sp_inst_1.INIT_RAM_3A = 256'h92CC31AC418C018C31CC32CE058CB2CC31AD280C92CD3C0092C0BBFF958DE40C;
defparam sp_inst_1.INIT_RAM_3B = 256'hE40C018D31AC32CD058CB2CC5D8DC00C018D31AC32CD058CB2CCB2CC058CB2CC;
defparam sp_inst_1.INIT_RAM_3C = 256'h058CB2CC8FFF01848ECC9BFF34040DAC280C8ECD24000000B7FF94043FFF958D;
defparam sp_inst_1.INIT_RAM_3D = 256'h72C4C076B076406300208063E076F0610184000CC59F018C31AC32CDB2CCB2CC;
defparam sp_inst_1.INIT_RAM_3E = 256'h098D280D72CC0D8D72CC818D31AC000C818D0D8C72CC0D8D0C0D72CCA2C0BEC0;
defparam sp_inst_1.INIT_RAM_3F = 256'h180D72CC058072CC0D8D72CC818DFD8C818C0D8C72CC058072CC018D140D72CC;

SP sp_inst_2 (
    .DO({sp_inst_2_dout_w[15:0],sp_inst_2_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_2}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_2.READ_MODE = 1'b0;
defparam sp_inst_2.WRITE_MODE = 2'b01;
defparam sp_inst_2.BIT_WIDTH = 16;
defparam sp_inst_2.BLK_SEL = 3'b001;
defparam sp_inst_2.RESET_MODE = "SYNC";
defparam sp_inst_2.INIT_RAM_00 = 256'hB2CC0000AECC00ACB2C48076707680630020C063B0760000BECC018C72CC098D;
defparam sp_inst_2.INIT_RAM_01 = 256'h0180100C40763076C0630020806370760000018DAECDB2CCF19F818C818C158C;
defparam sp_inst_2.INIT_RAM_02 = 256'h40763076C0630020406330760000018C100C40763076C0630020406330760000;
defparam sp_inst_2.INIT_RAM_03 = 256'h707680630020406330760000102C040C40763076C06300204063307600000420;
defparam sp_inst_2.INIT_RAM_04 = 256'h698072CC72C4C076B07640630020806370760000042C0DAC040CB2CDB2C48076;
defparam sp_inst_2.INIT_RAM_05 = 256'hA2CD318CD60CA2CC31ACB2CDB1ACFD8C1FEC018D218CD60CA2C0B2CCA18C72CC;
defparam sp_inst_2.INIT_RAM_06 = 256'hB5CDFC0D118CD60C018E118CD60C2400018D01AD118CD60C018D118CD60C018D;
defparam sp_inst_2.INIT_RAM_07 = 256'h0000BECC5D8C018C118CD10C7ECC008CC076B07640630020C063B0760000018D;
defparam sp_inst_2.INIT_RAM_08 = 256'hC076A076B06140630020C063B0760000018D7ECDD10CF1AC080C098D5D8CBECC;
defparam sp_inst_2.INIT_RAM_09 = 256'hBECC018C72CC72CC058C72CC73FF0184BECC7FFF34040DAC280CBECD300072C4;
defparam sp_inst_2.INIT_RAM_0A = 256'h42C752C662C572C4C076A076B06140630020C063A076B0610184000CC59FBECC;
defparam sp_inst_2.INIT_RAM_0B = 256'h92CD52CC5000B2C092CC72CC0C00F7FFB40492CC300C72CC1D8072CC258042CC;
defparam sp_inst_2.INIT_RAM_0C = 256'h058CB2CC92CC000709A035CC92CE52CDC1AC35CDC2CEB2CD5DCC00070980B1AE;
defparam sp_inst_2.INIT_RAM_0D = 256'hA2CC1D8DB2CCA2CD7400A2CC31CC358CB5CE31ADB2CEB2CD62CCB19F92CCB2CC;
defparam sp_inst_2.INIT_RAM_0E = 256'h82CC1400818CC18C818C82CC198D240C82CD82CC000C0800C18C31ACC2CDFD8C;
defparam sp_inst_2.INIT_RAM_0F = 256'h0020C063A076B0610184000C8C0CA2CCA2CCFD8CA2CC07FF0184818C5D8C818C;
defparam sp_inst_2.INIT_RAM_10 = 256'h62CC62CC918C82CC72CB62CA52C942C832C722C612C532C40076E076F0618063;
defparam sp_inst_2.INIT_RAM_11 = 256'h32CD058CB2CC92CC040CE5AC940C7ECD7ECC018C31AC32CDB2CC8000B2C0A2CC;
defparam sp_inst_2.INIT_RAM_12 = 256'hA2CC7BFF0184018CA2CC0180018C31AC518C00AC898DADAC4C0D6D8C018C31AC;
defparam sp_inst_2.INIT_RAM_13 = 256'h058CB2CCA2CC118CA2CCEFFF0184818C018CA2CC9800B2CC058CB2CCA2CC118C;
defparam sp_inst_2.INIT_RAM_14 = 256'h3000B2CC058CB2CCA2CC118CA2CC83FF018492C528060007018CA2CC6800B2CC;
defparam sp_inst_2.INIT_RAM_15 = 256'h018CA2CCF800B2CC058CB2CCA2CC118CA2CC4BFF018492C528060407018CA2CC;
defparam sp_inst_2.INIT_RAM_16 = 256'h08060007018CA2CCC000B2CC058CB2CCA2CC118CA2CC13FF018492C520060007;
defparam sp_inst_2.INIT_RAM_17 = 256'h018492C540060007018CA2CC8800B2CC058CB2CCA2CC118CA2CCDBFF018492C5;
defparam sp_inst_2.INIT_RAM_18 = 256'h058CB2CC3800B2CC058CB2CCB3FF94045000B2CC058CB2CCA2CC118CA2CCA3FF;
defparam sp_inst_2.INIT_RAM_19 = 256'h058CB2CC92CC31AC418C018C31CC32CE058CB2CC31AD280C92CD3C0092C0B2CC;
defparam sp_inst_2.INIT_RAM_1A = 256'hBBFF958DE40C018D31AC32CD058CB2CCD98DC00C018D31AC32CD058CB2CCB2CC;
defparam sp_inst_2.INIT_RAM_1B = 256'hB2CC058CB2CC92CC31AC418C018C31CC32CE058CB2CC31AD280C92CD3C0092C0;
defparam sp_inst_2.INIT_RAM_1C = 256'h94043FFF958DE40C018D31AC32CD058CB2CC5D8DC00C018D31AC32CD058CB2CC;
defparam sp_inst_2.INIT_RAM_1D = 256'hB5CC3C0DB2CE4D80B2CC6FFF01847ECC7BFF34040DAC280C7ECD2400000097FF;
defparam sp_inst_2.INIT_RAM_1E = 256'hB2CCE59F82CDFD8D82CC0000000000000000140082CCCD8C00AC3580000709A0;
defparam sp_inst_2.INIT_RAM_1F = 256'h80767076806300208063E076F0610184000C759F018C31AC32CDB2CCB2CC058C;
defparam sp_inst_2.INIT_RAM_20 = 256'h406330760000BD80400C40763076C0630020806370760184B2CCB2CC600CB2C0;
defparam sp_inst_2.INIT_RAM_21 = 256'hB2CCB2C480766076706180630020406330760000BD8C400C40763076C0630020;
defparam sp_inst_2.INIT_RAM_22 = 256'hC076A076B061406300208063607670610000018DB2CC008D6BFF1180B2CC0180;
defparam sp_inst_2.INIT_RAM_23 = 256'h280031AC018C72CC118D72CC1DAC018C72CC118D72CC118D72CC008D33FF72C4;
defparam sp_inst_2.INIT_RAM_24 = 256'hB06140630020C063A076B061018431AC118C72CC31ADB2CD018C72CCB2CCFC0C;
defparam sp_inst_2.INIT_RAM_25 = 256'hB2CDB2C43FFF018492CC140007FF018492CCCBFFA2C092C0B2C072C4C076A076;
defparam sp_inst_2.INIT_RAM_26 = 256'h01848D8CB2CCB2C480766076706180630020C063A076B0610000BFFFE9AC72CC;
defparam sp_inst_2.INIT_RAM_27 = 256'h018431AC018C002CB2CDB2C48076607670618063002080636076706100007BFF;
defparam sp_inst_2.INIT_RAM_28 = 256'h9FFF018431ACA00CB2CDB2C48076607670618063002080636076706100003BFF;
defparam sp_inst_2.INIT_RAM_29 = 256'h0D80018CB2CD058DB2CC2000A2C5B2C480767076806300208063607670610000;
defparam sp_inst_2.INIT_RAM_2A = 256'hA2CCA2CCFD8CA2CC018D018CB2CCCDAC018CA2CE058EA2CC018DB2CC4400000C;
defparam sp_inst_2.INIT_RAM_2B = 256'hB2CC018C318CD70CA2C0B2C072C4C076B0764063002080637076018431AC018C;
defparam sp_inst_2.INIT_RAM_2C = 256'h818D3D8C818C958CB2CC158D72CC818DFD8C818CA58CB2CCA2CC018C218CD70C;
defparam sp_inst_2.INIT_RAM_2D = 256'hA2CC098D72CC818D7D8C818CC18CA2CC0D8D72CC818D7D8C818CB2CC118D72CC;
defparam sp_inst_2.INIT_RAM_2E = 256'hC063B0760000018D72CC818DFD8C818C918CA2CC058D72CC818DFD8C818CA98C;
defparam sp_inst_2.INIT_RAM_2F = 256'hB2CC118D040DB2CC1180118CB2CC118D300C118DB2CCB2C48076707680630020;
defparam sp_inst_2.INIT_RAM_30 = 256'hB1AE600C098DB2CC018D000DD70C0D8D040DB2CC11800D8CB2CC118D7C0C0D8D;
defparam sp_inst_2.INIT_RAM_31 = 256'hF00C018EB2CC31ADA98C81EC00070980B1CFF00C058EB2CCC18D81CC00070980;
defparam sp_inst_2.INIT_RAM_32 = 256'h218CD70C358D81ED000709A0B5CF900D19AEB2CD31AC918C81EC00070980B1CF;
defparam sp_inst_2.INIT_RAM_33 = 256'h7D8C0D8CB2CC31AD958C81EC00070980B1CF340C118EB2CCA58D158CB2CC018D;
defparam sp_inst_2.INIT_RAM_34 = 256'h80766076706180630020806370760000018D000D118CD70C018D318CD70C31AD;
defparam sp_inst_2.INIT_RAM_35 = 256'h40630020806360767061000063FFA2C40C0083FFA2C41180BECCBECCA2C5008C;
defparam sp_inst_2.INIT_RAM_36 = 256'h31CCB2CC040E018DD60C318062CCB2CC72CC698D7C0C72CD62C572C4C076B076;
defparam sp_inst_2.INIT_RAM_37 = 256'h6800018D39ADD60C018E31CCB2CC040E018DD60C9000018DB9ADD60C018E300C;
defparam sp_inst_2.INIT_RAM_38 = 256'h2800418DB9ADD60C018E300C31CCB2CC040E418DD60C318062CCB2CC818C72CC;
defparam sp_inst_2.INIT_RAM_39 = 256'hC076B07640630020C063B0760000418D39ADD60C018E31CCB2CC040E418DD60C;
defparam sp_inst_2.INIT_RAM_3A = 256'h018E300C31CCB2CC040E118DD60C318062CCB2CC72CC698D7C0C72CD62C572C4;
defparam sp_inst_2.INIT_RAM_3B = 256'h818C72CC6800118D39ADD60C018E31CCB2CC040E118DD60C9000118DB9ADD60C;
defparam sp_inst_2.INIT_RAM_3C = 256'h518DD60C2800518DB9ADD60C018E300C31CCB2CC040E518DD60C318062CCB2CC;
defparam sp_inst_2.INIT_RAM_3D = 256'h018CD40C40763076C0630020C063B0760000518D39ADD60C018E31CCB2CC040E;
defparam sp_inst_2.INIT_RAM_3E = 256'h62CCB2C062C572C4C076B07640630020406330760000018D81AD11ADD40C818D;
defparam sp_inst_2.INIT_RAM_3F = 256'h118CD60C018E118CD60C018DB5CDFDADFFED118CD60C018E118CD60C4180318C;

SP sp_inst_3 (
    .DO({sp_inst_3_dout_w[15:0],sp_inst_3_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_3}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_3.READ_MODE = 1'b0;
defparam sp_inst_3.WRITE_MODE = 2'b01;
defparam sp_inst_3.BIT_WIDTH = 16;
defparam sp_inst_3.BLK_SEL = 3'b001;
defparam sp_inst_3.RESET_MODE = "SYNC";
defparam sp_inst_3.INIT_RAM_00 = 256'h72CC2000218D72CCB1AD300C018C62CC218D72CC2980118C62CC018D35CD000D;
defparam sp_inst_3.INIT_RAM_01 = 256'h62CC118D72CC018D72CC31AD018C62CC018D72CC218D72CC31AD018C62CC218D;
defparam sp_inst_3.INIT_RAM_02 = 256'h118D72CC31AD018C62CC118D72CC25AC040C218D62CC118D72CCB1AD300C018C;
defparam sp_inst_3.INIT_RAM_03 = 256'h318D72CC31AD018C62CC318D72CC118D72CCB1AD300C018C62CC118D72CC2400;
defparam sp_inst_3.INIT_RAM_04 = 256'h8076707680630020C063B0760000018D72CCB1AD300C018C62CC018D72CC2400;
defparam sp_inst_3.INIT_RAM_05 = 256'h806300208063707600003180B2CC218D040DB2CC118D040DB2CC0180B2CCB2C4;
defparam sp_inst_3.INIT_RAM_06 = 256'h707680630020806370760000318DB2CC31ADA2CC318DB2CCA2C5B2C480767076;
defparam sp_inst_3.INIT_RAM_07 = 256'h806370760000C18D35CDB2CDD60CC18E300CB2CCD18DA9ADB4ADD60CB2C48076;
defparam sp_inst_3.INIT_RAM_08 = 256'hC076A076B06140630020406330760000D18DA9ADB4ADD60C40763076C0630020;
defparam sp_inst_3.INIT_RAM_09 = 256'hB2CC000709A035CCA2CE018D62CC098D800D72CCA2CC018CF42CB2C062C572C4;
defparam sp_inst_3.INIT_RAM_0A = 256'h62CC118D62CC058D72CC818DA18CB2CC018D72CC818DB2CCB2CCFD8C898CB2CC;
defparam sp_inst_3.INIT_RAM_0B = 256'h72CC1180198C62CC098D72CC818D31AC000C818D31AC1D8C62CC818D31AC198C;
defparam sp_inst_3.INIT_RAM_0C = 256'h8076707680630020C063A076B06100003C00D2041D8D72CC158D62CC118D100D;
defparam sp_inst_3.INIT_RAM_0D = 256'h1D80B2CC198D080DB2CC158DA80DB2CC118D800DB2CC018D81AD030DB2CCB2C4;
defparam sp_inst_3.INIT_RAM_0E = 256'h818D018C818C118CB2CC2580A2CCA2C5B2C48076707680630020806370760000;
defparam sp_inst_3.INIT_RAM_0F = 256'h80630020806370760000118DB2CC818DB1ACFC0C818D118CB2CC2400118DB2CC;
defparam sp_inst_3.INIT_RAM_10 = 256'h70610000118D400DD20C0D8DAECDB2CC8400B2C4AECC00ACB2C4807660767061;
defparam sp_inst_3.INIT_RAM_11 = 256'h818C92CC818DA2CC3400B2C492C6A2C5B2C48076607670618063002080636076;
defparam sp_inst_3.INIT_RAM_12 = 256'hB2C4807660767061806300208063607670610000118DB2CC818D818C818C31AC;
defparam sp_inst_3.INIT_RAM_13 = 256'h108400A40185AECCAECC058CAECC2980AACCC800B2C4AACC01ACAECC00CD00AC;
defparam sp_inst_3.INIT_RAM_14 = 256'h400DD20C0D8DAECDB2CCA7FFE08400A40185AECCAECCB1ACF80CAECD2800CFFF;
defparam sp_inst_3.INIT_RAM_15 = 256'h118C72CC1000BECC118C72CC72C4C076B076406300208063607670610000118D;
defparam sp_inst_3.INIT_RAM_16 = 256'hBECCBECC118C72CC72C4C076B07640630020C063B0760000ED9F098CBECCBECC;
defparam sp_inst_3.INIT_RAM_17 = 256'hA076B06140630020C063B0760000118D72CC818D118C818C118C72CC2180118C;
defparam sp_inst_3.INIT_RAM_18 = 256'hBECCBECC818C818C818C9D8C7ACC7ACCFD8C7ACC76CC01AC7ACC00AD008CC076;
defparam sp_inst_3.INIT_RAM_19 = 256'h818C118CD20CEBFFD20447FFD20401850006BECC7BFF90840084018501A676CD;
defparam sp_inst_3.INIT_RAM_1A = 256'h0185818C7ACC1FFF1084008401857ACC7ACCFD8C7ACC3FFF4084008411805D8C;
defparam sp_inst_3.INIT_RAM_1B = 256'h03FFD204018576CCE3FFD084008411805D8C818C118CD20C8FFFD2043BFFD204;
defparam sp_inst_3.INIT_RAM_1C = 256'h000023FFD20463FFD2040405ABFFF084008411805D8C818C118CD20C57FFD204;
defparam sp_inst_3.INIT_RAM_1D = 256'h818C9D8C7ACC7ACCFD8C7ACC7ACC008CC076A076B06140630020C063A076B061;
defparam sp_inst_3.INIT_RAM_1E = 256'hD20CA3FFD204FFFFD20401850006BECC33FF908400840185BECCBECC818C818C;
defparam sp_inst_3.INIT_RAM_1F = 256'h7ACC7ACCFD8C7ACCE3FFF084008401857ACCF7FF1084008411805D8C818C118C;
defparam sp_inst_3.INIT_RAM_20 = 256'h0406BECC9BFFA084008411805D8C818C118CD20C47FFD204F3FFD2040185818C;
defparam sp_inst_3.INIT_RAM_21 = 256'hD204200500065FFFB084008411805D8C818C118CD20C0BFFD20467FFD2040185;
defparam sp_inst_3.INIT_RAM_22 = 256'hD80C8076707680630020C063A076B0610184BACCBACC0D8CD20CD3FFD204CFFF;
defparam sp_inst_3.INIT_RAM_23 = 256'h0000E9AC040CB2CDB2CC018C218CD80C1400B2CC018C218CD80C018D000D218C;
defparam sp_inst_3.INIT_RAM_24 = 256'h218CD80C1400B2CC018C218CD80C52C662C572C4C076B0764063002080637076;
defparam sp_inst_3.INIT_RAM_25 = 256'h52CD018D62CD118CD80C018DB5CDFDADFFED72CED80CE9AC040CB2CDB2CC018C;
defparam sp_inst_3.INIT_RAM_26 = 256'h80630020C063B0760000018D040D218CD80C1400018D0C0D218CD80C19AC040C;
defparam sp_inst_3.INIT_RAM_27 = 256'hB1CCFD8C01ECBD8E098CB2CC31ADC18C058CB2CCE18D018CB2CCB2C480767076;
defparam sp_inst_3.INIT_RAM_28 = 256'h0000018D218CD68C31AD3D8C118CB2CC31ADB1CC018C002CA18E0D8CB2CC31AD;
defparam sp_inst_3.INIT_RAM_29 = 256'h31ADB1CC800CD98E058CB2CCE18D018CB2CCB2C4807670768063002080637076;
defparam sp_inst_3.INIT_RAM_2A = 256'h318CD68C358D11ADB2CD31AC018CA18C0D8CB2CC31ADB1CC7E0CC18E098CB2CC;
defparam sp_inst_3.INIT_RAM_2B = 256'h01ECBD8E098CB2CCC18D018CB2CCB2C48076707680630020806370760000018D;
defparam sp_inst_3.INIT_RAM_2C = 256'h158CB2CC31AD018CAD8C118CB2CC31ADB1CC00ECB18E0D8CB2CC31ADB1CCFD8C;
defparam sp_inst_3.INIT_RAM_2D = 256'h058C218CB2CC31AD098C858C1D8CB2CC31ADFD8C918C198CB2CC31AD018CA18C;
defparam sp_inst_3.INIT_RAM_2E = 256'h018D118CD60C2580B2CCB2C48076707680630020806370760000018DD68C31AD;
defparam sp_inst_3.INIT_RAM_2F = 256'h806370760000018DB5CDFC0D118CD60C018E118CD60C2400018D01AD118CD60C;
defparam sp_inst_3.INIT_RAM_30 = 256'h818CFD8C818C018C31AC018CD68C018D898CBACCBACC008C8076707680630020;
defparam sp_inst_3.INIT_RAM_31 = 256'h018C31AC018CD68C018D898CBACCBACC008C8076707680630020806370760184;
defparam sp_inst_3.INIT_RAM_32 = 256'h0000018D09ADD68C018DD68C40763076C0630020806370760184818CFD8C818C;
defparam sp_inst_3.INIT_RAM_33 = 256'h80630020406330760000018D05ADD68C018DD68C40763076C063002040633076;
defparam sp_inst_3.INIT_RAM_34 = 256'hBACDFD8C018C31AC018CD68C018D898CBECCBACC01ACBECC00AD008C80767076;
defparam sp_inst_3.INIT_RAM_35 = 256'h70768063002080637076000001AC398C35ED01ADD68D01AF89ADBECD01AEE1AD;
defparam sp_inst_3.INIT_RAM_36 = 256'h018C31AC018CD68C018D898CBECC018EE18CBACCBACC01ACBECC00AD008C8076;
defparam sp_inst_3.INIT_RAM_37 = 256'hA076B0614063002080637076000001AC31CC35ED01ADD68D01AF89ADBECDFD8C;
defparam sp_inst_3.INIT_RAM_38 = 256'h2C0CBACDBACC058CBACC53FF018401A57ECD818CBACC2800BAC07ECC008CC076;
defparam sp_inst_3.INIT_RAM_39 = 256'hA6CC400CA2CC400C3ECC008C0076E076F06100630020C063A076B0610000D58D;
defparam sp_inst_3.INIT_RAM_3A = 256'h8ECC200C8ACC200C86C082CC0C0C1FFF0184A2CCB2CC040CAECC040CAACC040C;
defparam sp_inst_3.INIT_RAM_3B = 256'h6ACC0C0C66CC0C0C62C05ECC0C0C5ACC040C52CCFC0C7FFF018482CC92CCFC0C;
defparam sp_inst_3.INIT_RAM_3C = 256'h63FF0404C3FF01843ECCF59F058C018CD68C0000BBFFC7FF018452CC72C06EC0;
defparam sp_inst_3.INIT_RAM_3D = 256'h008CDBFF0184818CB2CC3C00B2C0407620763061C06300200063E076F0610000;
defparam sp_inst_3.INIT_RAM_3E = 256'hB2C017FF10840084C18D2C0CB2CDB2CC058CB2CC218D31CCC2CE898CB2CC018D;
defparam sp_inst_3.INIT_RAM_3F = 256'hC98D2C0CB2CDB2CC058CB2CCEBFFD08400840185218C31ACC2CD898CB2CC3400;

SP sp_inst_4 (
    .DO({sp_inst_4_dout_w[15:0],sp_inst_4_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_4}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_4.READ_MODE = 1'b0;
defparam sp_inst_4.WRITE_MODE = 2'b01;
defparam sp_inst_4.BIT_WIDTH = 16;
defparam sp_inst_4.BLK_SEL = 3'b001;
defparam sp_inst_4.RESET_MODE = "SYNC";
defparam sp_inst_4.INIT_RAM_00 = 256'h00204063207630610000A7FF708400840185AECCAECC3D8C818C018C118CD68C;
defparam sp_inst_4.INIT_RAM_01 = 256'h318CDA0C018D11ADB2CD218CDA0C0180118CDA0C0180DA0CB2C4807670768063;
defparam sp_inst_4.INIT_RAM_02 = 256'h818D018CD40C2180518CB2CC018D35CDDA0C518DB2CC018EDA0C018D21ADB2CD;
defparam sp_inst_4.INIT_RAM_03 = 256'hDA0C618DB2CC018EDA0C018D35CDDA0C418DB2CC018EDA0C018D81AD05ADD40C;
defparam sp_inst_4.INIT_RAM_04 = 256'h040DB2CC018D01ADF42DB2CCB2C48076707680630020806370760000018D35CD;
defparam sp_inst_4.INIT_RAM_05 = 256'hB2CC218D01AD026DB2CC118DFDAD002DB2CC418D100DB2CC518D080DB2CC618D;
defparam sp_inst_4.INIT_RAM_06 = 256'h018D05ADDA0C018DDA0C1D80B2CCB2C480767076806300208063707600003180;
defparam sp_inst_4.INIT_RAM_07 = 256'h3980B2CCB2C48076707680630020806370760000018DF9ADDA0C018DDA0C1800;
defparam sp_inst_4.INIT_RAM_08 = 256'hDA0C018DDA0C3800018D81AD05ADD40C818D018CD40C018D09ADDA0C018DDA0C;
defparam sp_inst_4.INIT_RAM_09 = 256'hB07640630020806370760000018D81ADB5CDF80DD40C818E018CD40C018DF5AD;
defparam sp_inst_4.INIT_RAM_0A = 256'hC063B0760184B2CCB2C00800B2CC040C1180B1AC72CC018DDA0CB2C072C4C076;
defparam sp_inst_4.INIT_RAM_0B = 256'hD40C818D018C0D8CD40C018D35CDB2CDDA0C018EDA0CB2C48076707680630020;
defparam sp_inst_4.INIT_RAM_0C = 256'h707601840000A2C5B2C48076707680630020806370760000018D81AD05AD0D8C;
defparam sp_inst_4.INIT_RAM_0D = 256'h0084AC0091AC080C72CD15AC040C72CD62C572C4C076A076B061406300208063;
defparam sp_inst_4.INIT_RAM_0E = 256'h2084008401C50186018C31AC918CB2CCE1AD008D058EB2CC4400B2C04BFFD084;
defparam sp_inst_4.INIT_RAM_0F = 256'h959F008C63FF508400840185018C31AC918CB2CC01AD008DB2CC058CB2CC0FFF;
defparam sp_inst_4.INIT_RAM_10 = 256'h008C1FFFA2C40185018C31AC918CB2CCE1AD008DA000B2C0A2CC118C62CC3800;
defparam sp_inst_4.INIT_RAM_11 = 256'hB2CC71AD008D218F31AC918CB2CCD1AD008D018E31AC918CB2CC31AD008D6980;
defparam sp_inst_4.INIT_RAM_12 = 256'hB2CC71AD008DB2CC058CB2CC40002FFFD084008401C501E60187318C31AC918C;
defparam sp_inst_4.INIT_RAM_13 = 256'h0185018C31AC918CB2CCB1AD008D399F008C7FFFC08400840185018C31AC918C;
defparam sp_inst_4.INIT_RAM_14 = 256'h0184000C00000800A3FF508400841400B3FF108400842580008C4FFF00840084;
defparam sp_inst_4.INIT_RAM_15 = 256'hB2CC1D8C38EC018D140D118CD10C33FF0076E076F06100630020C063A076B061;
defparam sp_inst_4.INIT_RAM_16 = 256'h1400A2CCCD8C00AC57FFC0840084E59FB2CDFD8DB2CC00000000000000001400;
defparam sp_inst_4.INIT_RAM_17 = 256'h00AC0BFFC084008442C542CCE18C008CE59FA2CDFD8DA2CC0000000000000000;
defparam sp_inst_4.INIT_RAM_18 = 256'h0084100532CC058C868CE59F92CDFD8D92CC0000000000000000140092CCCD8C;
defparam sp_inst_4.INIT_RAM_19 = 256'h22CC200CE59F82CDFD8D82CC0000000000000000140082CCCD8C00ACBFFFC084;
defparam sp_inst_4.INIT_RAM_1A = 256'h72CDFD8D72CC0000000000000000140072CCCD8C00AC73FFC0840084018522CC;
defparam sp_inst_4.INIT_RAM_1B = 256'h0000000000000000140062CC918C1C6C93FFA7FF50040405B3FF04040405E59F;
defparam sp_inst_4.INIT_RAM_1C = 256'h52CC0000000000000000140052CC918C1C6C5FFF04040405E59F62CDFD8D62CC;
defparam sp_inst_4.INIT_RAM_1D = 256'h40630020406330760184000C40763076C0638BFF23FF04040005E59F52CDFD8D;
defparam sp_inst_4.INIT_RAM_1E = 256'hC000040C1BFF60840084198D0C0C72CD118D040C72CD62C572C4C076A076B061;
defparam sp_inst_4.INIT_RAM_1F = 256'h0184018C218C62CC2000A2CC040C11AC080C72CD92C4FC000184018C118C62CC;
defparam sp_inst_4.INIT_RAM_20 = 256'hB2CD97FFD0840084018531AC92CCB2CD21801D8CB2CC5C00B2C0A2CC008CCC00;
defparam sp_inst_4.INIT_RAM_21 = 256'h0184000CA1ACA2CCB2CDB2CC058CB2CC73FF708400840185818C018C31AC92CC;
defparam sp_inst_4.INIT_RAM_22 = 256'h198D0C0C72CD118D040C72CD62C572C4C076A076B06140630020C063A076B061;
defparam sp_inst_4.INIT_RAM_23 = 256'hA2CC040C11AC080C72CD92C4E8000184018C118C62CCCC00040C07FFE0840084;
defparam sp_inst_4.INIT_RAM_24 = 256'h018D898CB2CC29800D8CB2CC6800B2C0A2CC008CB8000184018C218C62CC2000;
defparam sp_inst_4.INIT_RAM_25 = 256'h53FFB08400840185018C31AC92CC018D898CB2CC7BFF20840084018531AC92CC;
defparam sp_inst_4.INIT_RAM_26 = 256'hC076A076B06140630020C063A076B0610184000C95ACA2CCB2CDB2CC058CB2CC;
defparam sp_inst_4.INIT_RAM_27 = 256'hB2C4D4000184018C118C62CC4800040CF3FF5084008419AC0C0C72CD62C572C4;
defparam sp_inst_4.INIT_RAM_28 = 256'h0020C063A076B0610184000C018DAECDB2CCAECC008CBC000184018C218C62CC;
defparam sp_inst_4.INIT_RAM_29 = 256'h118C62CC4400040C63FF9084008419AC0C0C72CD62C572C4C076A076B0614063;
defparam sp_inst_4.INIT_RAM_2A = 256'hB0610184000C018DA2CDB2CCA2C42C000184018C218C62CCB2C444000184018C;
defparam sp_inst_4.INIT_RAM_2B = 256'h018D058C72CC41ACC00C018D72CCB2C072C4C076A076B06140630020C063A076;
defparam sp_inst_4.INIT_RAM_2C = 256'h19ACC00C018D72CC3400A2CC400C92CC080C19AC600C018D058C72CC19ACE00C;
defparam sp_inst_4.INIT_RAM_2D = 256'h280CA2CD82CC018C31AC92CC72CD5400A2CC280C92C06400A2CC200C92CC040C;
defparam sp_inst_4.INIT_RAM_2E = 256'hA2CCB2CD258DE40C82CD318DBC0C82CD0C00C5AC200CA2CD15AC400CA2CDDDAC;
defparam sp_inst_4.INIT_RAM_2F = 256'h82CC31ADA2CCB2CD258D980C82CD318D800C82CD8400B2CC418C31AC82CC31AD;
defparam sp_inst_4.INIT_RAM_30 = 256'h258C31AC82CC31ADA2CCB2CD258D180C82CD318D000C82CD4C00B2CCA58C31AC;
defparam sp_inst_4.INIT_RAM_31 = 256'hA2CCB2CD25AC82CDC18CA2CC358DBC0C82CD500054007FFF808400841400B2CC;
defparam sp_inst_4.INIT_RAM_32 = 256'h31AC92CC72CD92CC058C92CC00002FFFA08400841000B2CC418C31AC82CC31AD;
defparam sp_inst_4.INIT_RAM_33 = 256'h0C0C72CD62C572C4C076A076B06140630020C063A076B0610184B2CCA19F018C;
defparam sp_inst_4.INIT_RAM_34 = 256'h0184018C218C62CCB2C4A7FF0184018C118C62CC6400040CC3FF4084008419AC;
defparam sp_inst_4.INIT_RAM_35 = 256'hB0610184000C5FFF90840084ABFFB2C4A2C504067BFF908400846BFFA2C48FFF;
defparam sp_inst_4.INIT_RAM_36 = 256'h13FFF08400640185018CD68C2BFF2084008480766076706180630020C063A076;
defparam sp_inst_4.INIT_RAM_37 = 256'hD0840064DBFFB08400640185018C318CD68CF7FFD08400640185018C218CD68C;
defparam sp_inst_4.INIT_RAM_38 = 256'h31CC018CD68C018E898CB2CC018D31AC018CD68C018D898CB2CC6000B2C0CFFF;
defparam sp_inst_4.INIT_RAM_39 = 256'h70610184000C9D8D2C0CB2CDB2CC058CB2CC77FFF0840064B2C501A60187018C;
defparam sp_inst_4.INIT_RAM_3A = 256'hB2CC3400B2C01FFF108400642BFF208400648076607670618063002080636076;
defparam sp_inst_4.INIT_RAM_3B = 256'h10840064C98D2C0CB2CDB2CC058CB2CCF3FF808400640185008C3FFF0184818C;
defparam sp_inst_4.INIT_RAM_3C = 256'hB2CDB2CC058CB2CCA3FF408400640185008C3BFF0184818CB2CC3400B2C0CFFF;
defparam sp_inst_4.INIT_RAM_3D = 256'h118C62CC62C572C4C076A076B061406300208063607670610184000CC98D2C0C;
defparam sp_inst_4.INIT_RAM_3E = 256'h00644800040C1FFF9084006419AC0C0C72CD5D80008CC7FFF08400640185018C;
defparam sp_inst_4.INIT_RAM_3F = 256'h018C118C62CC0C006FFF0184BACCBACC008CF7FF0184018C218C62CC0BFFA084;

SP sp_inst_5 (
    .DO({sp_inst_5_dout_w[15:0],sp_inst_5_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_5}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_5.READ_MODE = 1'b0;
defparam sp_inst_5.WRITE_MODE = 2'b01;
defparam sp_inst_5.BIT_WIDTH = 16;
defparam sp_inst_5.BLK_SEL = 3'b001;
defparam sp_inst_5.RESET_MODE = "SYNC";
defparam sp_inst_5.INIT_RAM_00 = 256'h108400641D80818CB1AC818C058C098C72CC818D058C008C4BFFC08400640185;
defparam sp_inst_5.INIT_RAM_01 = 256'h53FF80840064C580008CEFFFB08400640185018C118C62CCB0000FFF8BFF8FFF;
defparam sp_inst_5.INIT_RAM_02 = 256'h018401A5BECCB6CD2400BEC03DAC0C0C72CDB6CC008C3FFF0184018C218C62CC;
defparam sp_inst_5.INIT_RAM_03 = 256'hD3FF0184018C318C62CC39AC100C72CD2000D98D2C0CBECDBECC058CBECC3FFF;
defparam sp_inst_5.INIT_RAM_04 = 256'h018C118C62CCD000040CA7FF10840064E000E7FF018401A5BECCB6CDBECC008C;
defparam sp_inst_5.INIT_RAM_05 = 256'h608400641980818CB1AC818C058C098C72CC818D058C008C0BFF108400640185;
defparam sp_inst_5.INIT_RAM_06 = 256'h058C098C72CC818D058C008CB3FF108400640185018C118C62CC74001BFF4FFF;
defparam sp_inst_5.INIT_RAM_07 = 256'h000C0800040CDFFF40840064EBFF308400642400BBFFBFFF1180818CB1AC818C;
defparam sp_inst_5.INIT_RAM_08 = 256'h0C0CF2CD9BFF60840064E2C5F2C4407620763061C0630020C063A076B0610184;
defparam sp_inst_5.INIT_RAM_09 = 256'hB2C457FF0184018C118CE2CC9C00040C73FF308400649BFF00044FFF0004298D;
defparam sp_inst_5.INIT_RAM_0A = 256'hB2CC63FF018422CC92C427FF0184018C318CE2CCA2C43FFF0184018C218CE2CC;
defparam sp_inst_5.INIT_RAM_0B = 256'h000C4BFF018422CC42CC31AC018CF42C92CD32CC31ACFD8C002CA2CD62CC898C;
defparam sp_inst_5.INIT_RAM_0C = 256'h72CD97FF7084006472C562C572C4C076A076B061406300204063207630610184;
defparam sp_inst_5.INIT_RAM_0D = 256'h458CB2CDB2C45FFF0184018C118C62CC3800040C7BFF808400646FFF1D8D040C;
defparam sp_inst_5.INIT_RAM_0E = 256'h62C572C4C076A076B06140630020C063A076B0610184000C6FFF018431ACE18C;
defparam sp_inst_5.INIT_RAM_0F = 256'h218C62CCB2C4DFFF0184018C118C62CCBC00040CFBFFE0840064198D080C72CD;
defparam sp_inst_5.INIT_RAM_10 = 256'h080CB2CD60009FFF20840064A2C583FFA2C421AC040CB2CDA2C4C7FF0184018C;
defparam sp_inst_5.INIT_RAM_11 = 256'h20840064A2C5ABFFA2C421AC0C0CB2CD380077FFA0840064A2C593FFA2C421AC;
defparam sp_inst_5.INIT_RAM_12 = 256'h72C4C076A076B06140630020C063A076B0610184000C3FFFF084006410004FFF;
defparam sp_inst_5.INIT_RAM_13 = 256'h2C00040CDBFF0084006443FF0004218D040C72CD9BFFFFFF0084006472C562C5;
defparam sp_inst_5.INIT_RAM_14 = 256'h80630020C063A076B0610184000CC7FF0FFFB2C4B2C4BFFF0184018C118C62CC;
defparam sp_inst_5.INIT_RAM_15 = 256'h0C00FC0C5BFF60840064198DE40CBECD118DBC0CBECDBECC008C807660767061;
defparam sp_inst_5.INIT_RAM_16 = 256'hA084006462C572C4C0769077A076B0614063002080636076706101843D8CBECC;
defparam sp_inst_5.INIT_RAM_17 = 256'h01A5E2CD018C118C62CC12CC02CDF2CEE2CF318C218D118E018F618C006C0FFF;
defparam sp_inst_5.INIT_RAM_18 = 256'h93FF808400649FFF10840064ABFF90840064B7FF508400643D80008C53FF0184;
defparam sp_inst_5.INIT_RAM_19 = 256'h6084006419AC100C72CDA180008CF7FF018401A5F2CD018C118C62CC6000000C;
defparam sp_inst_5.INIT_RAM_1A = 256'h31B7280C008D8FFF0184018CB2CCA2CC318C62CCB2CC218C62CC1C00040C4FFF;
defparam sp_inst_5.INIT_RAM_1B = 256'h31B7280C008D4FFF0184018C0D8CB2CC92CC32EC008C6FFF0184018C058CB2CC;
defparam sp_inst_5.INIT_RAM_1C = 256'h31B7280C008D0FFF0184018C198CB2CC82CC32EC008C2FFF0184018C118CB2CC;
defparam sp_inst_5.INIT_RAM_1D = 256'hA2CC31B7280C008DD3FF0184018CA2CC72CC32EC008CEFFF0184018C1D8CB2CC;
defparam sp_inst_5.INIT_RAM_1E = 256'hA2CC31B7280C008D93FF0184018C0D8CA2CC62CC32EC008CB3FF0184018C058C;
defparam sp_inst_5.INIT_RAM_1F = 256'hA2CC31B7280C008D53FF0184018C198CA2CC52CC32EC008C73FF0184018C118C;
defparam sp_inst_5.INIT_RAM_20 = 256'h72CC498D7C0C72CD558082CC5D8D300C82CD42CC32EC008C33FF0184018C1D8C;
defparam sp_inst_5.INIT_RAM_21 = 256'h0D8DF00C42CD118DF00C52CD1D8D600C62CD298D740C72CD11AC080C82CD4180;
defparam sp_inst_5.INIT_RAM_22 = 256'h818C52CCC2CC818C42CCFC00040C2FFF30840064198032CC32CC000C0800040C;
defparam sp_inst_5.INIT_RAM_23 = 256'h00040185C2CCD6CC818C92CCD2CC818C82CCCECC818C72CCCACC818C62CCC6CC;
defparam sp_inst_5.INIT_RAM_24 = 256'h6084006419AC100C72CD4980008C37FF018401A502CD018C118C62CCA00033FF;
defparam sp_inst_5.INIT_RAM_25 = 256'h31B7280C008DCFFF0184018C22CC12CC318C62CC22CC218C62CC5C00040C8FFF;
defparam sp_inst_5.INIT_RAM_26 = 256'h31B7280C008D8FFF0184018C0D8C22CC02CC32EC008CAFFF0184018C058C22CC;
defparam sp_inst_5.INIT_RAM_27 = 256'h12CC31B7280C008D53FF0184018C12CCF2CC32EC008C6FFF0184018C118C22CC;
defparam sp_inst_5.INIT_RAM_28 = 256'h12CC31B7280C008D13FF0184018C0D8C12CCE2CC32EC008C33FF0184018C058C;
defparam sp_inst_5.INIT_RAM_29 = 256'h12CC31B7280C008DD3FF0184018C198C12CCD2CC32EC008CF3FF0184018C118C;
defparam sp_inst_5.INIT_RAM_2A = 256'hF2CC498D7C0CF2CD558002CC5D8D300C02CDC2CC32EC008CB3FF0184018C1D8C;
defparam sp_inst_5.INIT_RAM_2B = 256'h0D8DF00CC2CD118DF00CD2CD1D8D600CE2CD298D740CF2CD11AC080C02CD4180;
defparam sp_inst_5.INIT_RAM_2C = 256'h818CD2CCA2CC818CC2CC7C00040CAFFF308400641980B2CCB2CC000C0800040C;
defparam sp_inst_5.INIT_RAM_2D = 256'h12CD018C118C62CC3800000CB2CC818C02CCAECC818CF2CCAACC818CE2CCA6CC;
defparam sp_inst_5.INIT_RAM_2E = 256'h818DB1ACC18C00ECA2CDA2C42BFF0184018C218C62CC8980008CCFFF018401A5;
defparam sp_inst_5.INIT_RAM_2F = 256'h918CA2CCB000040CE3FF408400641980818C31AC818C058CB1CC458C018CA2CE;
defparam sp_inst_5.INIT_RAM_30 = 256'hF7FF0404018582CCA3FFC084006411AC040C72CD9000000C82CC3D8CA2CC92CC;
defparam sp_inst_5.INIT_RAM_31 = 256'h006472C562C652C722CC82CC32CC86CC42CC8ACC52CC8ECC62CC92CC72CC96CC;
defparam sp_inst_5.INIT_RAM_32 = 256'h40630020C0639077A076B0610184000C33FFA084006442C532C622C74BFFB084;
defparam sp_inst_5.INIT_RAM_33 = 256'hD3FF6084006417FF1D8D040C72CDEFFF5084006472C562C572C4C076A076B061;
defparam sp_inst_5.INIT_RAM_34 = 256'h0020C063A076B0610184000C97FFB2C4B2C4B7FF0184018C118C62CC2800040C;
defparam sp_inst_5.INIT_RAM_35 = 256'hB06101840000C3FFD2040185A2CCD7FF0184A2CC62C572C4C076A076B0614063;
defparam sp_inst_5.INIT_RAM_36 = 256'h040C17FFC084006419AC100C72CD62C572C4C076A076B06140630020C063A076;
defparam sp_inst_5.INIT_RAM_37 = 256'hD3FF0184018C218C62CCBECC008CEFFF0184018C118C62CC03FF70840064C400;
defparam sp_inst_5.INIT_RAM_38 = 256'h598C31AC598CBACC598D9D8CBECCB6CC008CB7FF0184018C318C62CCBACC008C;
defparam sp_inst_5.INIT_RAM_39 = 256'h7BFF018401A5AACCB6CD67FFE08400640185AACC7BFF008400640185B6CCAACC;
defparam sp_inst_5.INIT_RAM_3A = 256'h006419AC0C0C72CD62C572C4C076A076B06140630020C063A076B0610184000C;
defparam sp_inst_5.INIT_RAM_3B = 256'hA2C4D7FF0184018C218C62CCB2C4EFFF0184018C118C62CC9800040C0BFFA084;
defparam sp_inst_5.INIT_RAM_3C = 256'h01849ACC9ACC31AC818CFD8C818CA2CC818DB1AC018C00EC818D9D8C818CB2CC;
defparam sp_inst_5.INIT_RAM_3D = 256'hF06100630020C063A076B0610184000C73FFD0840064018596CC96CC008C13FF;
defparam sp_inst_5.INIT_RAM_3E = 256'hA2C417FF0184018C218C22CCB2C42FFF0184018C118C22CC22C532C40076E076;
defparam sp_inst_5.INIT_RAM_3F = 256'h92CC000C0800040C0D8D100C32CD118D080C32CD1D8D080CA2CD298D1C0CB2CD;

SP sp_inst_6 (
    .DO({sp_inst_6_dout_w[15:0],sp_inst_6_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_6}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_6.READ_MODE = 1'b0;
defparam sp_inst_6.WRITE_MODE = 2'b01;
defparam sp_inst_6.BIT_WIDTH = 16;
defparam sp_inst_6.BLK_SEL = 3'b001;
defparam sp_inst_6.RESET_MODE = "SYNC";
defparam sp_inst_6.INIT_RAM_00 = 256'h006497FF20840064A3FFE0840064318092CC72CC008CBFFF0184018C318C22CC;
defparam sp_inst_6.INIT_RAM_01 = 256'h018D35CDB2CDB18CD60C918EA2CC7800018D010D118CD60CBC00040C8BFF6084;
defparam sp_inst_6.INIT_RAM_02 = 256'h0185B18C31AC580C82CD82CC018CC18CD60C018D01ADB18CD60C018DB18CD60C;
defparam sp_inst_6.INIT_RAM_03 = 256'hB5CDFDADFEED118CD60C018E118CD60C899F72CC72CCFD8C72CC07FFA0840064;
defparam sp_inst_6.INIT_RAM_04 = 256'h19AC080C72CD62C572C4C076A076B061406300200063E076F0610184000C018D;
defparam sp_inst_6.INIT_RAM_05 = 256'hD60C018ED60C1D80B2CCB2C46BFF0184018C118C62CC2800040C87FFE0840064;
defparam sp_inst_6.INIT_RAM_06 = 256'hD60CAC0061AC080CB2CD1580B2CC3DAC040CB2CDBD8D080CB2CD018D35CD040D;
defparam sp_inst_6.INIT_RAM_07 = 256'h018ED60C018DB5CDFDADFFEDD60C018ED60C8C00018DB5CDFDADFFEDD60C018E;
defparam sp_inst_6.INIT_RAM_08 = 256'h000DD60C018ED60C018DB5CDFDADFFEDD60C018ED60C5400018D35CD000DD60C;
defparam sp_inst_6.INIT_RAM_09 = 256'hB0610184000C018D000D118CD60C1800040C77FF6084006418000000018D35CD;
defparam sp_inst_6.INIT_RAM_0A = 256'hCC0C018DFC0D218CCC0C018DFC0D118CCC0C80766076706180630020C063A076;
defparam sp_inst_6.INIT_RAM_0B = 256'h00640FFF018D35CD000DCC0CB1AEFD8C07ECB2CDB000B2CC000C018D400D618C;
defparam sp_inst_6.INIT_RAM_0C = 256'hA2CC018D01ADA2CC018D31AC000CA2CD2C00A2CCB2CC018D000DCC0CCBFF0084;
defparam sp_inst_6.INIT_RAM_0D = 256'h018CB2CC018D35CD000DCC0CB1AEFD8C07ECB2CDCD8DA2CDFD8CB2CCA2CC118C;
defparam sp_inst_6.INIT_RAM_0E = 256'h018C31CC000CA2CE018DA2CC3800A2CCB2CC6000B2CC000C4DAC040CB2CDB2CC;
defparam sp_inst_6.INIT_RAM_0F = 256'h040CB2CDB2CC018CB2CCC18DA2CDFD8CB2CCA2CC118CA2CC03FFF084004411AC;
defparam sp_inst_6.INIT_RAM_10 = 256'h19AC080C72CD62C572C4C076A076B061406300208063607670610184000C9DAC;
defparam sp_inst_6.INIT_RAM_11 = 256'hF7FFD10411AC040CB2CDB2C46BFF0184018C118C62CC6400040C87FF30840044;
defparam sp_inst_6.INIT_RAM_12 = 256'hA076B0610184000C0800040C2BFFC08400441800DFFFD18411AC080CB2CD3000;
defparam sp_inst_6.INIT_RAM_13 = 256'h008C93FF118D800DCE0C018D480DCE0C62C572C4C076A076B06140630020C063;
defparam sp_inst_6.INIT_RAM_14 = 256'h0076E076F06100630020C063A076B06101840000BBFF608400440185BACCBACC;
defparam sp_inst_6.INIT_RAM_15 = 256'h92C457FF0184018C118C22CCE800040C73FF7084004419AC080C32CD22C532C4;
defparam sp_inst_6.INIT_RAM_16 = 256'h31ADB2CC82CD4000B2C082CCA18CA2CC9400A2C072CC000C43FF2084004482C0;
defparam sp_inst_6.INIT_RAM_17 = 256'h0044BD8DFC0CB2CDB2CC058CB2CC018D81AD01CD31ACB2CC62CD018E31AC000C;
defparam sp_inst_6.INIT_RAM_18 = 256'h004469AC72CCA2CDA2CC058CA2CC63FF018462C5000631AC82CC92CDCBFF8084;
defparam sp_inst_6.INIT_RAM_19 = 256'h080C32CD22C532C40076E076F061006300200063E076F0610184000C8BFF9084;
defparam sp_inst_6.INIT_RAM_1A = 256'h13FF2084004482C092C427FF0184018C118C22CC2800040C43FF8084004419AC;
defparam sp_inst_6.INIT_RAM_1B = 256'h8000B2C033FF018462C5000631AC82CC92CD82CCA18CA2CCD400A2C072CC000C;
defparam sp_inst_6.INIT_RAM_1C = 256'h018C31ACB2CC62CD45AC818C018C31CC000C31CEB2CC82CE018D31ACB2CC62CD;
defparam sp_inst_6.INIT_RAM_1D = 256'hB2CDB2CC058CB2CC1C0067FFB084004401C5018631AC000C31ADB2CC82CD018E;
defparam sp_inst_6.INIT_RAM_1E = 256'h0184000C1BFFD084004429AC72CCA2CDA2CC058CA2CC3FFF508400447D8DFC0C;
defparam sp_inst_6.INIT_RAM_1F = 256'hD3FFE084004419AC080C72CD62C572C4C076A076B061406300200063E076F061;
defparam sp_inst_6.INIT_RAM_20 = 256'h31AC020CB2CDC3FFB2C4A7FFA0840044B2C4B7FF0184018C118C62CC4800040C;
defparam sp_inst_6.INIT_RAM_21 = 256'h82C092C022C532C40076E076F06100630020C063A076B0610184000CAFFF0184;
defparam sp_inst_6.INIT_RAM_22 = 256'h37FF92C41BFFE084004401857ACC7ACC008CF3FF118D800DCE0C018D480DCE0C;
defparam sp_inst_6.INIT_RAM_23 = 256'hB2C082CCA18CA2CC9400A2C062CC000CF3FF1084004423FF018431AC020C92CD;
defparam sp_inst_6.INIT_RAM_24 = 256'hB2CC058CB2CC018D81AD01CD31ACB2CC52CD018E31AC000C31ADB2CC82CD4000;
defparam sp_inst_6.INIT_RAM_25 = 256'hA2CC058CA2CC5FFFD08400441FFF018452C5000631AC82CC92CDBD8DFC0CB2CD;
defparam sp_inst_6.INIT_RAM_26 = 256'h82CCA18CA2CCD400A2C062CC000C2FFF808400443BFF7084004469AC62CCA2CD;
defparam sp_inst_6.INIT_RAM_27 = 256'h31CEB2CC82CE018D31ACB2CC52CD8000B2C04FFF018452C5000631AC82CC92CD;
defparam sp_inst_6.INIT_RAM_28 = 256'h018631AC000C31ADB2CC82CD018E018C31ACB2CC52CD45AC818C018C31CC000C;
defparam sp_inst_6.INIT_RAM_29 = 256'h058CA2CC5BFFC08400447D8DFC0CB2CDB2CC058CB2CC1C0083FF2084004401C5;
defparam sp_inst_6.INIT_RAM_2A = 256'h60767061806300200063E076F0610184000C37FFF084004429AC62CCA2CDA2CC;
defparam sp_inst_6.INIT_RAM_2B = 256'h098C100C43FF018482CC47FF6184D60C200500065BFF4184D60C080500068076;
defparam sp_inst_6.INIT_RAM_2C = 256'h60767061018400007BFF8184D60C018582CCB2CC040CA2CC040C92CC040C82CC;
defparam sp_inst_6.INIT_RAM_2D = 256'h406300208063607670610184000C57FFA2C5B2C4807660767061806300208063;
defparam sp_inst_6.INIT_RAM_2E = 256'h62C572C4C076A076B06140630020C063B0760184000CB2C062C572C4C076B076;
defparam sp_inst_6.INIT_RAM_2F = 256'hB2C0DDAC004CB2CDB2CC118CB2CC018031AC000CB2CD2000B2C007FF70840044;
defparam sp_inst_6.INIT_RAM_30 = 256'h004CB2CDB2CC118CB2CC01AC01CC018D31AC000CB2CD018E31AC020CB2CD3800;
defparam sp_inst_6.INIT_RAM_31 = 256'h018E31AC000CB2CD3DAC018C31CC020CB2CE018D31AC000CB2CD6C00B2C0C5AC;
defparam sp_inst_6.INIT_RAM_32 = 256'h91AC004CB2CDB2CC118CB2CC2BFF50840044B2C501C60187018C31AC020CB2CD;
defparam sp_inst_6.INIT_RAM_33 = 256'h00445C05C0C60046407620763061C0630020C063A076B0610184000C0180000C;
defparam sp_inst_6.INIT_RAM_34 = 256'h0046407620763061C063002040632076306100006BFF8184D60C0405CBFF3084;
defparam sp_inst_6.INIT_RAM_35 = 256'h3061C063002040632076306100001FFF8184D60C08057FFF008400447005F0C6;
defparam sp_inst_6.INIT_RAM_36 = 256'h4063207630610000D3FF8184D60C100533FFD0840044840520C6004640762076;
defparam sp_inst_6.INIT_RAM_37 = 256'h000087FF8184D60C2005E7FFA0840044980550C60046407620763061C0630020;
defparam sp_inst_6.INIT_RAM_38 = 256'hD60C40059BFF70840044AC0580C60046407620763061C0630020406320763061;
defparam sp_inst_6.INIT_RAM_39 = 256'h40840044C005B0C60046407620763061C063002040632076306100003BFF8184;
defparam sp_inst_6.INIT_RAM_3A = 256'hE0C60046407620763061C06300204063207630610000EFFF8184D60C80054FFF;
defparam sp_inst_6.INIT_RAM_3B = 256'h20763061C06300204063207630610000A3FF8184D60C000503FF10840044D405;
defparam sp_inst_6.INIT_RAM_3C = 256'h0020406320763061000057FF8184D60C0005B7FFE0840044EC0510C600464076;
defparam sp_inst_6.INIT_RAM_3D = 256'h306100000BFF8184D60C00056BFFB0840044000540C60046407620763061C063;
defparam sp_inst_6.INIT_RAM_3E = 256'h8184D60C00051FFF80840044180570C60046407620763061C063002040632076;
defparam sp_inst_6.INIT_RAM_3F = 256'hD3FF508400443005A0C60046407620763061C06300204063207630610000BFFF;

SP sp_inst_7 (
    .DO({sp_inst_7_dout_w[15:0],sp_inst_7_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_7}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_7.READ_MODE = 1'b0;
defparam sp_inst_7.WRITE_MODE = 2'b01;
defparam sp_inst_7.BIT_WIDTH = 16;
defparam sp_inst_7.BLK_SEL = 3'b001;
defparam sp_inst_7.RESET_MODE = "SYNC";
defparam sp_inst_7.INIT_RAM_00 = 256'h4805D0C60046407620763061C0630020406320763061000073FF8184D60C0005;
defparam sp_inst_7.INIT_RAM_01 = 256'h407620763061C0630020406320763061000027FF8184D60C000587FF20840044;
defparam sp_inst_7.INIT_RAM_02 = 256'hC06300204063207630610000DBFF8184D60C00253BFFF08400445C0500C60046;
defparam sp_inst_7.INIT_RAM_03 = 256'h2076306100008FFF8184D60C0045EFFFC0840044700530C60046407620763061;
defparam sp_inst_7.INIT_RAM_04 = 256'h43FF8184D60C0085A3FF90840044880560C60046407620763061C06300204063;
defparam sp_inst_7.INIT_RAM_05 = 256'h010557FF60840044A00590C60046407620763061C06300204063207630610000;
defparam sp_inst_7.INIT_RAM_06 = 256'h0044BC05C0C60046407620763061C06300204063207630610000F7FF8184D60C;
defparam sp_inst_7.INIT_RAM_07 = 256'h0046407620763061C06300204063207630610000ABFF8184D60C02050BFF3084;
defparam sp_inst_7.INIT_RAM_08 = 256'h3061C063002040632076306100005FFF8184D60C0405BFFF00840044D405F0C6;
defparam sp_inst_7.INIT_RAM_09 = 256'h406320763061000013FF8184D60C080573FFD0840044EC0520C6004640762076;
defparam sp_inst_7.INIT_RAM_0A = 256'h0000C7FF8184D60C100527FFA0840044040550C60046407620763061C0630020;
defparam sp_inst_7.INIT_RAM_0B = 256'hD60C2005DBFF708400441C0580C60046407620763061C0630020406320763061;
defparam sp_inst_7.INIT_RAM_0C = 256'h408400443005B0C60046407620763061C063002040632076306100007BFF8184;
defparam sp_inst_7.INIT_RAM_0D = 256'hE0C60046407620763061C063002040632076306100002FFF8184D60C40058FFF;
defparam sp_inst_7.INIT_RAM_0E = 256'h20763061C06300204063207630610000E3FF8184D60C800543FF108400444405;
defparam sp_inst_7.INIT_RAM_0F = 256'h0020406320763061000097FF8184D60C0005F7FFE08400445C0510C600464076;
defparam sp_inst_7.INIT_RAM_10 = 256'h306100004BFF8184D60C0005ABFFB0840044740540C60046407620763061C063;
defparam sp_inst_7.INIT_RAM_11 = 256'h8184D60C00055FFF808400448C0570C60046407620763061C063002040632076;
defparam sp_inst_7.INIT_RAM_12 = 256'h13FF50840044A405A0C60046407620763061C06300204063207630610000FFFF;
defparam sp_inst_7.INIT_RAM_13 = 256'hBC05D0C60046407620763061C06300204063207630610000B3FF8184D60C0005;
defparam sp_inst_7.INIT_RAM_14 = 256'h407620763061C0630020406320763061000067FF8184D60C0005C7FF20840044;
defparam sp_inst_7.INIT_RAM_15 = 256'hC063002040632076306100001BFF8184D60C00057BFFF0840024D40500C60046;
defparam sp_inst_7.INIT_RAM_16 = 256'h207630610000CFFF8184D60C00052FFFC0840024F00530C60046407620763061;
defparam sp_inst_7.INIT_RAM_17 = 256'h83FF8184D60C0005E3FF90840024080560C60046407620763061C06300204063;
defparam sp_inst_7.INIT_RAM_18 = 256'h000597FF60840024200590C60046407620763061C06300204063207630610000;
defparam sp_inst_7.INIT_RAM_19 = 256'h018D000DF18CD60C80766076706180630020406320763061000037FF8184D60C;
defparam sp_inst_7.INIT_RAM_1A = 256'h92CCA2CD92CC018C818CD60CA2CC318C818CD60C3BFFF0840024D00580C60046;
defparam sp_inst_7.INIT_RAM_1B = 256'h018C31AC898CB2CCD1AD002D2180058CB1ACB2CCA2CD4000B2C00000A2CCB1AC;
defparam sp_inst_7.INIT_RAM_1C = 256'h807660767061806300208063607670610000BD8D7C0CB2CDB2CC058CB2CC0181;
defparam sp_inst_7.INIT_RAM_1D = 256'h7061806300208063607670610000A7FFB2CC018C118CD60C018D020DF18CD60C;
defparam sp_inst_7.INIT_RAM_1E = 256'hD60CB6CC3D8C818C018C118CD68CBACCFD8C818CC18C018C118CD68C80766076;
defparam sp_inst_7.INIT_RAM_1F = 256'h8063607670610000E3FFB08400240185BACC018D3C0D118CD68C018D040DF18C;
defparam sp_inst_7.INIT_RAM_20 = 256'h0020806370760000BECC018C098CD18C018D080DF18CD60C8076707680630020;
defparam sp_inst_7.INIT_RAM_21 = 256'hF00DF18CD60C018E118CD60CB2CC7D8CCD8C018C118CD60C8076607670618063;
defparam sp_inst_7.INIT_RAM_22 = 256'hD60C17FF008400240180018C31AC018C002C898DB2CC718D400CB2CD018DB5CD;
defparam sp_inst_7.INIT_RAM_23 = 256'h0800018DB5CDFDADFEED118CD60C018E118CD60CFBFF308400243C000180118C;
defparam sp_inst_7.INIT_RAM_24 = 256'h058C9ECC9ECC018C158CD40C8076607670618063002080636076706100000000;
defparam sp_inst_7.INIT_RAM_25 = 256'h218CFF0C018D518CFF0C018D818C058C018CB18CFF0C4980008C33FF00045980;
defparam sp_inst_7.INIT_RAM_26 = 256'hD10C6C00BECC018C118CD10CA2C09180118C9ECC33FF0004EBFF50040185018C;
defparam sp_inst_7.INIT_RAM_27 = 256'h280DD10CA2C01980A2CC2C00A2CC040C018D340DD10C1DAC340C82CD82CC018C;
defparam sp_inst_7.INIT_RAM_28 = 256'hD40C1580218C9ECC919F058CBECCBECC018C118CD10C018D82CDD10C1000018D;
defparam sp_inst_7.INIT_RAM_29 = 256'h407620763061C06300208063607670610000018DFC0D0D8CD40C018D200D0D8C;
defparam sp_inst_7.INIT_RAM_2A = 256'h0000000000000000000000000020406320763061000027FF43FFE084002457FF;
defparam sp_inst_7.INIT_RAM_2B = 256'h1F081F081F081F081F081F081F081F081DEC0066636238373433300070756177;
defparam sp_inst_7.INIT_RAM_2C = 256'h1F081F081F081F081E8C1E8C1E8C1E8C1E8C1E8C1E8C1E8C1E8C1E041F081F08;
defparam sp_inst_7.INIT_RAM_2D = 256'h1F081F081F081F081F081F081F081F081F081F081F081F081F081F081F081F08;
defparam sp_inst_7.INIT_RAM_2E = 256'h1F081F081F081F081F081F081F081F081F081F081F081F081F081F081F081F08;
defparam sp_inst_7.INIT_RAM_2F = 256'h1F081F081F081F081F081F081F081F081F081D0C1CA41D7C1F081F081F081F08;
defparam sp_inst_7.INIT_RAM_30 = 256'h273C273C273C273C26201DB41F081F081CD41F081C781F081F081DB41D441F08;
defparam sp_inst_7.INIT_RAM_31 = 256'h26C026C026C026C026C026C026C026C026C02638273C273C273C273C273C273C;
defparam sp_inst_7.INIT_RAM_32 = 256'h273C273C273C273C273C273C273C273C273C273C273C273C273C273C273C273C;
defparam sp_inst_7.INIT_RAM_33 = 256'h273C273C273C273C273C273C273C273C273C273C273C273C273C273C273C273C;
defparam sp_inst_7.INIT_RAM_34 = 256'h273C273C273C273C273C254024D825B0273C273C273C273C273C273C273C273C;
defparam sp_inst_7.INIT_RAM_35 = 256'h0A0D25E8273C273C2508273C24AC273C273C25E82578273C273C273C273C273C;
defparam sp_inst_7.INIT_RAM_36 = 256'h72645F6576650A0D0A0D30252072612061720A0D000078327830646465766365;
defparam sp_inst_7.INIT_RAM_37 = 256'h61650A0D78253D7261570A0D2D2D63616E2D2D2D000025783D2061642C202578;
defparam sp_inst_7.INIT_RAM_38 = 256'h0A0D6E770A0D000A250978253D7261520A206120200A20787830646465636544;
defparam sp_inst_7.INIT_RAM_39 = 256'h310909383730300909343330300909300A0D564F6E750A0D6E77696C0A0D0000;
defparam sp_inst_7.INIT_RAM_3A = 256'h2D2D6156430A0000250900002509000056620A0D00002509006C65730A0D3131;
defparam sp_inst_7.INIT_RAM_3B = 256'h2D2D005D756E3E72613C645B316400005D74655B00007865007830207079654B;
defparam sp_inst_7.INIT_RAM_3C = 256'h6568726F73736464706D2D2D005D756E3E72613C645B3464747973736464706D;
defparam sp_inst_7.INIT_RAM_3D = 256'h2D2D3E6561763E72613C6D5B316D747320642D2D0000646E6D6F2070685B0000;
defparam sp_inst_7.INIT_RAM_3E = 256'h77206572612069642D2D3E6561763E72613C6D5B346D00656220657261206964;
defparam sp_inst_7.INIT_RAM_3F = 256'h616C000073657265745B000070686863745B00686F7400002D2D765B00760064;

SP sp_inst_8 (
    .DO({sp_inst_8_dout_w[15:0],sp_inst_8_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_8}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_8.READ_MODE = 1'b0;
defparam sp_inst_8.WRITE_MODE = 2'b01;
defparam sp_inst_8.BIT_WIDTH = 16;
defparam sp_inst_8.BLK_SEL = 3'b001;
defparam sp_inst_8.RESET_MODE = "SYNC";
defparam sp_inst_8.INIT_RAM_00 = 256'h7565775B70756177000073657961645B00796564005D6574656D2065635B656D;
defparam sp_inst_8.INIT_RAM_01 = 256'h65722070695B000032695D747420775B64775D747420725B00006164005D6574;
defparam sp_inst_8.INIT_RAM_02 = 256'h64773E7261673C20646469682077695B00003269656C736520632D2D005D6C61;
defparam sp_inst_8.INIT_RAM_03 = 256'h646120632D2D3E7261673C20646469682072695B00003269746920632D2D3E61;
defparam sp_inst_8.INIT_RAM_04 = 256'h6873665F735B00006F6300006E3C6564625B7465616200632D2D005D615B6461;
defparam sp_inst_8.INIT_RAM_05 = 256'h2074755B0074697500003C2064742D2D5D79635B006D695F6F63005D616C6E69;
defparam sp_inst_8.INIT_RAM_06 = 256'h6574775F735B000070736573655F735B736170735D74695F735B746970737469;
defparam sp_inst_8.INIT_RAM_07 = 256'h00745D69655B0000695F70676873665F735B687366735D64725F735B00007073;
defparam sp_inst_8.INIT_RAM_08 = 256'h7F287F1448907F107EFC7EE8477C7EE47EE07ED843207ED05D4C4E5B0000554E;
defparam sp_inst_8.INIT_RAM_09 = 256'h7FCC7FC84CE07FC47FAC7F984A407F947F7C7F6849B07F647F587F4443487F3C;
defparam sp_inst_8.INIT_RAM_0A = 256'h7FCC802053A880187FCC800453147FFC7FCC7FEC52147FE47FCC7FDC4F607FD4;
defparam sp_inst_8.INIT_RAM_0B = 256'h808880745D40806C7FCC80605CBC805C7FCC8050559C80487FCC803854AC8030;
defparam sp_inst_8.INIT_RAM_0C = 256'h7FCC811C611C8114810C81045F78810080F480D85E9880D080C480A05D8C8098;
defparam sp_inst_8.INIT_RAM_0D = 256'h7FCC818C64C881847FCC8178641C8170816081586BA8814C7FCC8134628C812C;
defparam sp_inst_8.INIT_RAM_0E = 256'h7FCC81DC686081D47FCC81C8666081C07FCC81B4653081AC7FCC81A067D08198;
defparam sp_inst_8.INIT_RAM_0F = 256'h00003A73616D630A82008208475C82007FCC81F46B7C81FC7FCC81F46B4881E8;
defparam sp_inst_8.INIT_RAM_10 = 256'h6761200A000A21646D6D2065666575204F52090A73252509090A0D0A3A642009;
defparam sp_inst_8.INIT_RAM_11 = 256'h203D756E0A0D203D656C0D733D207473000042410A0D240A0D0A6D6320706820;
defparam sp_inst_8.INIT_RAM_12 = 256'h6761200A20782520093A3025200A00003E6D3C2072643C2064206761200A0A0D;
defparam sp_inst_8.INIT_RAM_13 = 256'h61763E72613C6D206761200A2078252000093830300A0D0A756E3E72613C6420;
defparam sp_inst_8.INIT_RAM_14 = 256'h0A2E7265756E656861676C6900003E6561763E72613C6D206761200A00003E65;
defparam sp_inst_8.INIT_RAM_15 = 256'h6574612064205056000D6D75203E646176206761200A0A2E7265756E61676C69;
defparam sp_inst_8.INIT_RAM_16 = 256'h30202020727453540A3A736E540A000A652065746120642050560A2074727320;
defparam sp_inst_8.INIT_RAM_17 = 256'h202072746E6820202020783830206D696C6F5354783830202020637353547838;
defparam sp_inst_8.INIT_RAM_18 = 256'h302032302031202020202020200A7838302020787830205D255B000065524320;
defparam sp_inst_8.INIT_RAM_19 = 256'h630A000025206C61616200003120303120392020202030203630203520202020;
defparam sp_inst_8.INIT_RAM_1A = 256'h200A0000637300006E496375200A3E686E773C206E696375200A00006E696176;
defparam sp_inst_8.INIT_RAM_1B = 256'h68633E686E773C206F646375200A68546F446375200A00006F64000063536375;
defparam sp_inst_8.INIT_RAM_1C = 256'h6567550A2E7272457570200A00006873002E6F506375200A00006F700000656E;
defparam sp_inst_8.INIT_RAM_1D = 256'h203E6E6E633C6874776F206E6420756F202020200920745F6F64746920686F74;
defparam sp_inst_8.INIT_RAM_1E = 256'h6863742020200A096C6C20686F742020200A206E7320756F2020202020202020;
defparam sp_inst_8.INIT_RAM_1F = 256'h6174203E646F65707465203A61730A0D00002E2E72612072697465700A0D6F68;
defparam sp_inst_8.INIT_RAM_20 = 256'h20726974203A61730A0D642567722E2E726120726974726F0A0D3E633C206D5F;
defparam sp_inst_8.INIT_RAM_21 = 256'h736D0A0D73750A0D3E6C3C203A336D3A73753A656D3C616C203A61730A0D6365;
defparam sp_inst_8.INIT_RAM_22 = 256'h3C20656B203A61730A0D000A3A63612E2E74747355206157656D0A0D00730A0D;
defparam sp_inst_8.INIT_RAM_23 = 256'h0000202E6974616C6964742061640A0D0A0D65626E20206561726E6F0A0D3E63;
defparam sp_inst_8.INIT_RAM_24 = 256'h6D3A20646D6D2D20616400002E657420732020736D6D68202D6D79792D206164;
defparam sp_inst_8.INIT_RAM_25 = 256'h732020726574206E7963716520746E697A482D20616400002E742074206F7373;
defparam sp_inst_8.INIT_RAM_26 = 256'h6220756F0A0D006D6170696C6E69000A65746172206B686300002E6563737020;
defparam sp_inst_8.INIT_RAM_27 = 256'h3025002030253230643230320D6573756F662D2061640D7A3836332020656C63;
defparam sp_inst_8.INIT_RAM_28 = 256'h2E2E6174747320670A0D8A188A148A108A0C662D692D732D682D64323A64253A;
defparam sp_inst_8.INIT_RAM_29 = 256'h61673C2064646968207769206761200A63652067203A61730A0D0000253A7261;
defparam sp_inst_8.INIT_RAM_2A = 256'h6572726470693C7269206761200A0078303D646178253D6164773E6164773E72;
defparam sp_inst_8.INIT_RAM_2B = 256'h3A6C0A0D003E6D69203E643C6C6520430A0D000A3230302061640A0D000A6464;
defparam sp_inst_8.INIT_RAM_2C = 256'h293128563129202C4F523428563029332C5052562820495F4129202C5F432930;
defparam sp_inst_8.INIT_RAM_2D = 256'h6761200A00647461636C0A0D6420202C203A3A760A0D636D6164282065723628;
defparam sp_inst_8.INIT_RAM_2E = 256'h002E0072656D61706E6F0A0D314F47202C305047202C5F4320306E3C65646220;
defparam sp_inst_8.INIT_RAM_2F = 256'h746973206761200A0D78303D0A0D0A202F31746975206761200A726F65206F63;
defparam sp_inst_8.INIT_RAM_30 = 256'h200A203E6461646173206761200A000A202E0A7474737469200A00003E72613C;
defparam sp_inst_8.INIT_RAM_31 = 256'h613C736173206761200A7825646420786174722072726B63630A000A61746461;
defparam sp_inst_8.INIT_RAM_32 = 256'h63650A0D656E206D676F0A0D0A747473617272700A7474737361200A00003E72;
defparam sp_inst_8.INIT_RAM_33 = 256'h2C78726F65206F630A0D61746D6179700A0D000A6F6463650A0D000A61747475;
defparam sp_inst_8.INIT_RAM_34 = 256'h544E54462E2E2E2E2E2E2E0A00003E2073256E756425656E20200A0D0000252C;
defparam sp_inst_8.INIT_RAM_35 = 256'h2E2E2E2E2E2E2E0A000A7830656E68434B3A49686F742D0A0D0A2E2E2E2E2E2E;
defparam sp_inst_8.INIT_RAM_36 = 256'h6F43000D2E2E2E2E2E2E2E432E2E2E2E2E2E2E0A0D0A2E2E2E2E2E2E4C495F54;
defparam sp_inst_8.INIT_RAM_37 = 256'h6F406EF46EA86E5C6E106DC46D786D2C6CE0000A747072656920656C72655420;
defparam sp_inst_8.INIT_RAM_38 = 256'h740073B47368731C72D07284723871EC71A07154710870BC707070246FD86F8C;
defparam sp_inst_8.INIT_RAM_39 = 256'h790079007900790079007900790078B07900761475C8757C753074E47498744C;
defparam sp_inst_8.INIT_RAM_3A = 256'h675F7865656C61687269616F675F786578CC7900790079007900790079007900;
defparam sp_inst_8.INIT_RAM_3B = 256'h656C61687269616F675F7865656C61687269616F675F7865656C61687269616F;
defparam sp_inst_8.INIT_RAM_3C = 256'h7269616F675F7865656C61687269616F675F7865656C61687269616F675F7865;
defparam sp_inst_8.INIT_RAM_3D = 256'h675F7865656C61687269626F675F7865656C61687269616F675F7865656C6168;
defparam sp_inst_8.INIT_RAM_3E = 256'h656C61687269626F675F7865656C61687269626F675F7865656C61687269626F;
defparam sp_inst_8.INIT_RAM_3F = 256'h7269626F675F7865656C61687269626F675F7865656C61687269626F675F7865;

SP sp_inst_9 (
    .DO({sp_inst_9_dout_w[15:0],sp_inst_9_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_9}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_9.READ_MODE = 1'b0;
defparam sp_inst_9.WRITE_MODE = 2'b01;
defparam sp_inst_9.BIT_WIDTH = 16;
defparam sp_inst_9.BLK_SEL = 3'b001;
defparam sp_inst_9.RESET_MODE = "SYNC";
defparam sp_inst_9.INIT_RAM_00 = 256'h675F7865656C61687269636F675F7865656C61687269626F675F7865656C6168;
defparam sp_inst_9.INIT_RAM_01 = 256'h656C61687269636F675F7865656C61687269636F675F7865656C61687269636F;
defparam sp_inst_9.INIT_RAM_02 = 256'h7269636F675F7865656C61687269636F675F7865656C61687269636F675F7865;
defparam sp_inst_9.INIT_RAM_03 = 256'h675F7865656C61687269646F675F7865656C61687269636F675F7865656C6168;
defparam sp_inst_9.INIT_RAM_04 = 256'h656C61687269646F675F7865656C61687269646F675F7865656C61687269646F;
defparam sp_inst_9.INIT_RAM_05 = 256'h7269646F675F7865656C61687269646F675F7865656C61687269646F675F7865;
defparam sp_inst_9.INIT_RAM_06 = 256'h000000007AC07AC90000656C61687865656C61687269646F675F7865656C6168;
defparam sp_inst_9.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_10 (
    .DO({sp_inst_10_dout_w[15:0],sp_inst_10_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_10}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_10.READ_MODE = 1'b0;
defparam sp_inst_10.WRITE_MODE = 2'b01;
defparam sp_inst_10.BIT_WIDTH = 16;
defparam sp_inst_10.BLK_SEL = 3'b001;
defparam sp_inst_10.RESET_MODE = "SYNC";
defparam sp_inst_10.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_11 (
    .DO({sp_inst_11_dout_w[15:0],sp_inst_11_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_11}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_11.READ_MODE = 1'b0;
defparam sp_inst_11.WRITE_MODE = 2'b01;
defparam sp_inst_11.BIT_WIDTH = 16;
defparam sp_inst_11.BLK_SEL = 3'b001;
defparam sp_inst_11.RESET_MODE = "SYNC";
defparam sp_inst_11.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_12 (
    .DO({sp_inst_12_dout_w[15:0],sp_inst_12_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_12}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_12.READ_MODE = 1'b0;
defparam sp_inst_12.WRITE_MODE = 2'b01;
defparam sp_inst_12.BIT_WIDTH = 16;
defparam sp_inst_12.BLK_SEL = 3'b001;
defparam sp_inst_12.RESET_MODE = "SYNC";
defparam sp_inst_12.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_13 (
    .DO({sp_inst_13_dout_w[15:0],sp_inst_13_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_13}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_13.READ_MODE = 1'b0;
defparam sp_inst_13.WRITE_MODE = 2'b01;
defparam sp_inst_13.BIT_WIDTH = 16;
defparam sp_inst_13.BLK_SEL = 3'b001;
defparam sp_inst_13.RESET_MODE = "SYNC";
defparam sp_inst_13.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_14 (
    .DO({sp_inst_14_dout_w[15:0],sp_inst_14_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_14}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_14.READ_MODE = 1'b0;
defparam sp_inst_14.WRITE_MODE = 2'b01;
defparam sp_inst_14.BIT_WIDTH = 16;
defparam sp_inst_14.BLK_SEL = 3'b001;
defparam sp_inst_14.RESET_MODE = "SYNC";
defparam sp_inst_14.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_15 (
    .DO({sp_inst_15_dout_w[15:0],sp_inst_15_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_15}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_15.READ_MODE = 1'b0;
defparam sp_inst_15.WRITE_MODE = 2'b01;
defparam sp_inst_15.BIT_WIDTH = 16;
defparam sp_inst_15.BLK_SEL = 3'b001;
defparam sp_inst_15.RESET_MODE = "SYNC";
defparam sp_inst_15.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_16 (
    .DO({sp_inst_16_dout_w[15:0],sp_inst_16_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_16.READ_MODE = 1'b0;
defparam sp_inst_16.WRITE_MODE = 2'b01;
defparam sp_inst_16.BIT_WIDTH = 16;
defparam sp_inst_16.BLK_SEL = 3'b001;
defparam sp_inst_16.RESET_MODE = "SYNC";
defparam sp_inst_16.INIT_RAM_00 = 256'h15005FFF00100380150003801500028029800010288000100386143850000015;
defparam sp_inst_16.INIT_RAM_01 = 256'h03BF15FF040003BF140004000015040014385FFF028029805800038015000380;
defparam sp_inst_16.INIT_RAM_02 = 256'h00000000000000004C0006484C00544403BD1500040003800406038814EC0406;
defparam sp_inst_16.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_17 (
    .DO({sp_inst_17_dout_w[15:0],sp_inst_17_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_1}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_17.READ_MODE = 1'b0;
defparam sp_inst_17.WRITE_MODE = 2'b01;
defparam sp_inst_17.BIT_WIDTH = 16;
defparam sp_inst_17.BLK_SEL = 3'b001;
defparam sp_inst_17.RESET_MODE = "SYNC";
defparam sp_inst_17.INIT_RAM_00 = 256'h29BE29BE29BE29BE29BE29BF29BF29BF29BF29BF29BF29BF29BF29BF15000400;
defparam sp_inst_17.INIT_RAM_01 = 256'h440003404400034044000340440003404000036E040029BE29BE29BE29BE29BE;
defparam sp_inst_17.INIT_RAM_02 = 256'h5000546950005465500054675000546750005466500054664400036044000342;
defparam sp_inst_17.INIT_RAM_03 = 256'h28BE28BE28BF28BF28BF28BF28BF28BF28BF28BF28BF15005000546840000341;
defparam sp_inst_17.INIT_RAM_04 = 256'h2900157F43FF03402A00157F0648040028BE28BE28BE28BE28BE28BE28BE28BE;
defparam sp_inst_17.INIT_RAM_05 = 256'h57FF03802A00001000170014580003800380038015E028BA1CC8298002BF4C00;
defparam sp_inst_17.INIT_RAM_06 = 256'h43FF03402A00157F58002A0000154C000280288057FF038053FF02BF02BF0044;
defparam sp_inst_17.INIT_RAM_07 = 256'h29BF29BF29BF29BF29BF150004004C0043FF03412A00157F53FF02802900157F;
defparam sp_inst_17.INIT_RAM_08 = 256'h29BE29BE29BE29BE29BE29BF29BF29BF29BF29BF29BF29BF29BF29BF29BF29BF;
defparam sp_inst_17.INIT_RAM_09 = 256'h03402880157F387229BE0400028029BE29BE29BE29BE29BE29BE29BE29BE29BE;
defparam sp_inst_17.INIT_RAM_0A = 256'h28BF28BF28BF28BF28BF28BF28BF28BF28BF150057FF28B51CC80648298043FF;
defparam sp_inst_17.INIT_RAM_0B = 256'h28BE28BE28BE28BE28BE28BE28BE28BE28BE28BF28BF28BF28BF28BF28BF28BF;
defparam sp_inst_17.INIT_RAM_0C = 256'h001529BF0280298002BF4C00040004000380040028BE28BE28BE28BE28BE28BE;
defparam sp_inst_17.INIT_RAM_0D = 256'h2A3F4000034000182A3F2A7F5000293F29BF288028BF29BF29BF29BF297F29BF;
defparam sp_inst_17.INIT_RAM_0E = 256'h001528BF001728BF28BF29BF001428BF001428BF29BF001728BF028029BF0040;
defparam sp_inst_17.INIT_RAM_0F = 256'h298002BF4C00028028800340298028BF28BF6FFF02802A3F293F02802A3F29BF;
defparam sp_inst_17.INIT_RAM_10 = 256'h28BF28BF29BF028028BF29002A00157F001028BF28BF500029BF29BF29BF0280;
defparam sp_inst_17.INIT_RAM_11 = 256'h290000672A00001028BF28BF157F500029BF43FF034000672A00157F03406BFF;
defparam sp_inst_17.INIT_RAM_12 = 256'h28BF157F47FF034000672A00157F03406BFF28BF001502BF28BF29BF028028BF;
defparam sp_inst_17.INIT_RAM_13 = 256'h29BF29BF29BF0280298002BF4C00028028800340290000672A00001028BF02BF;
defparam sp_inst_17.INIT_RAM_14 = 256'h0340500029BF6FFF028028BF29BF028028BF29002A00157F001028BF28BF5000;
defparam sp_inst_17.INIT_RAM_15 = 256'h157F001028BF28BF290000672A00001028BF28BF157F47FF034000672A00157F;
defparam sp_inst_17.INIT_RAM_16 = 256'h00672A00157F034050006BFF28BF28BF29BF028028BF29BF028028BF29002A00;
defparam sp_inst_17.INIT_RAM_17 = 256'h03406BFF28BF28BF29BF028028BF290000672A00001028BF28BF157F47FF0340;
defparam sp_inst_17.INIT_RAM_18 = 256'h00672A00157F290000670380157F00672A00157F0280298002BF4C0002802880;
defparam sp_inst_17.INIT_RAM_19 = 256'h157F00672A00157F0280298002BF4C0002802880034029000067001402BF157F;
defparam sp_inst_17.INIT_RAM_1A = 256'h298002BF4C00028028800340290000670380157F00672A00157F290000670380;
defparam sp_inst_17.INIT_RAM_1B = 256'h02802880288000152A3F57FF57FD0015028002BF57FF293F028029BF02802980;
defparam sp_inst_17.INIT_RAM_1C = 256'h02BF4C00028028802880034047FF0340001557FF034002802980298002BF4C00;
defparam sp_inst_17.INIT_RAM_1D = 256'h28802880034057FE57FC0015028002BF57FE57FF293F028029BF028029802980;
defparam sp_inst_17.INIT_RAM_1E = 256'h57FC0015028002BF57FE293F293F293F293F02BE02802980298002BF4C000280;
defparam sp_inst_17.INIT_RAM_1F = 256'h02802980298002BF4C0002802880288000152A4002BF57FE57FC0015028002BF;
defparam sp_inst_17.INIT_RAM_20 = 256'h29BF004428BF293F006728BF29BF004428BF293F006728BF293F02BF29BF29BF;
defparam sp_inst_17.INIT_RAM_21 = 256'h4C00028028802880034057FE57FE57FB0015028002BF57FD57FE293F006728BF;
defparam sp_inst_17.INIT_RAM_22 = 256'h29BF004428BF293F006728BF293F028029BF29BF29BF29BF02802980298002BF;
defparam sp_inst_17.INIT_RAM_23 = 256'h28BF57FB0015028002BF57FD57FE293F006728BF29BF004428BF293F006728BF;
defparam sp_inst_17.INIT_RAM_24 = 256'h29BF29BF29BF02802980298002BF4C00028028802880034057FD57FD57FB28BF;
defparam sp_inst_17.INIT_RAM_25 = 256'h28BF29BF004428BF293F006728BF29BF004428BF293F006728BF293F028029BF;
defparam sp_inst_17.INIT_RAM_26 = 256'h4C00028028802880034057FC57FB28BF28BF57FA0015028002BF57FC293F0067;
defparam sp_inst_17.INIT_RAM_27 = 256'h02BE4C0002802880288003405406157F00152A3F293F001502802980298002BF;
defparam sp_inst_17.INIT_RAM_28 = 256'h57FF028029BF001128BE640028BE400028BE29BE29BE29BE29BE028129812981;
defparam sp_inst_17.INIT_RAM_29 = 256'h28BE293E001002BF28BF0000002A5C00002128BF28BE500029BF29BF28BE5000;
defparam sp_inst_17.INIT_RAM_2A = 256'h00130013001228BF28BF28BE47FF28BF29BF028028BF29BF002A5C00002128BF;
defparam sp_inst_17.INIT_RAM_2B = 256'h028028BF29BF00155000283E001002BF02BF28BF600028BF28BF500029BF0015;
defparam sp_inst_17.INIT_RAM_2C = 256'h28BF29BF02BF28BF57FE001500670281006728BF500000670280006728BF6000;
defparam sp_inst_17.INIT_RAM_2D = 256'h5C000280283F500029BF02802980298002BF4C000281288128810015001563FF;
defparam sp_inst_17.INIT_RAM_2E = 256'h28800015001547FF283F293F2A0028BF29BF028028BF57FE00152A3F57FE0280;
defparam sp_inst_17.INIT_RAM_2F = 256'h0280298029802980298029802980298029BF02812980298002BE4C0002802880;
defparam sp_inst_17.INIT_RAM_30 = 256'h29BF02805C020280283F293F2A00001028BF28BF500329BF29BF28BF29BF02BF;
defparam sp_inst_17.INIT_RAM_31 = 256'h288028BF4C002880001002B91C0000406802028102BF2800001028BF028028BF;
defparam sp_inst_17.INIT_RAM_32 = 256'h028028BF57FD00150067288028BF500229BF028028BF29BF028028BF57FE0015;
defparam sp_inst_17.INIT_RAM_33 = 256'h28BF29BF028028BF57FD001528BF02800015288028BF500229BF028028BF29BF;
defparam sp_inst_17.INIT_RAM_34 = 256'h29BF028028BF29BF028028BF57FC001528BF02800280288028BF500229BF0280;
defparam sp_inst_17.INIT_RAM_35 = 256'h28BF500129BF028028BF29BF028028BF57FC001528BF02800015288028BF5001;
defparam sp_inst_17.INIT_RAM_36 = 256'h0015288028BF500129BF028028BF29BF028028BF57FC001528BF028000152880;
defparam sp_inst_17.INIT_RAM_37 = 256'h29BF028028BF57FB0280500129BF028028BF29BF028028BF57FC001528BF0280;
defparam sp_inst_17.INIT_RAM_38 = 256'h001002BF2800001028BF028028BF001C028028BF500029BF29BF028028BF5001;
defparam sp_inst_17.INIT_RAM_39 = 256'h2800001028BF028028BF67FD02802800001028BF028028BF29BF028028BF29BF;
defparam sp_inst_17.INIT_RAM_3A = 256'h29BF001002BF2800001028BF028028BF001C028028BF500029BF53FD67FF0280;
defparam sp_inst_17.INIT_RAM_3B = 256'h02802800001028BF028028BF67FD02802800001028BF028028BF29BF028028BF;
defparam sp_inst_17.INIT_RAM_3C = 256'h028028BF57FA00152A3F57FA02805C000280283F5000034057FA028053FD67FF;
defparam sp_inst_17.INIT_RAM_3D = 256'h29BF0280298002BF4C000281288028800015001547FC2800001028BF28BF29BF;
defparam sp_inst_17.INIT_RAM_3E = 256'h290002BF28BF290028BF0067001502BE00672A0028BF2900028028BF29BF293F;
defparam sp_inst_17.INIT_RAM_3F = 256'h028028BF290028BF290028BF0067034100672A0028BF290028BF2900028028BF;

SP sp_inst_18 (
    .DO({sp_inst_18_dout_w[15:0],sp_inst_18_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_2}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_18.READ_MODE = 1'b0;
defparam sp_inst_18.WRITE_MODE = 2'b01;
defparam sp_inst_18.BIT_WIDTH = 16;
defparam sp_inst_18.BLK_SEL = 3'b001;
defparam sp_inst_18.RESET_MODE = "SYNC";
defparam sp_inst_18.INIT_RAM_00 = 256'h28BF0340293F001529BF0280298002BF4C00028028800340293F2A0028BF2900;
defparam sp_inst_18.INIT_RAM_01 = 256'h040003800280298002BF4C0002802880034029002A3F28BF43FF034000672A00;
defparam sp_inst_18.INIT_RAM_02 = 256'h0280298002BF4C00028028800340040003800280298002BF4C00028028800340;
defparam sp_inst_18.INIT_RAM_03 = 256'h298002BF4C00028028800340040103800280298002BF4C000280288003400401;
defparam sp_inst_18.INIT_RAM_04 = 256'h400028BF29BF0280298002BF4C0002802880034004010380040128BF29BF0280;
defparam sp_inst_18.INIT_RAM_05 = 256'h28BF0380157F29BF001028BF001403BF140028800380157F29BF29BF004028BF;
defparam sp_inst_18.INIT_RAM_06 = 256'h001402B90380157F28800380157F5000298003860380157F28800380157F2980;
defparam sp_inst_18.INIT_RAM_07 = 256'h0340293F000028800380157F293F00150280298002BF4C000280288003402980;
defparam sp_inst_18.INIT_RAM_08 = 256'h02802980298002BF4C0002802880034029802A3F157F5BFF0280034000002A3F;
defparam sp_inst_18.INIT_RAM_09 = 256'h293F2A0028BF29BF028028BF57FF00152A3F57FF02805C000280283F500029BF;
defparam sp_inst_18.INIT_RAM_0A = 256'h29BE29BE29BE29BE02812981298102BE4C000280288028800015001547FF283F;
defparam sp_inst_18.INIT_RAM_0B = 256'h28BF28BE500029BF29BF28BE500057FE028029BF001128BE640028BE400028BE;
defparam sp_inst_18.INIT_RAM_0C = 256'h028028BF29BF002A5C00002128BF28BE293E001002BF28BF0000002A5C000021;
defparam sp_inst_18.INIT_RAM_0D = 256'h28BF600028BF28BF500029BF001500130013001228BF28BF28BE47FF28BF29BF;
defparam sp_inst_18.INIT_RAM_0E = 256'h28BF500000670280006728BF6000028028BF29BF00155000283E001002BF02BF;
defparam sp_inst_18.INIT_RAM_0F = 256'h4C000281288128810015001563FF28BF29BF02BF28BF57FE0015006702810067;
defparam sp_inst_18.INIT_RAM_10 = 256'h28BF29BF02BF0280298029802980298029802980298029BF02812980298002BE;
defparam sp_inst_18.INIT_RAM_11 = 256'h28BF028028BF29BF02805C020280283F293F2A00001028BF28BF500329BF29BF;
defparam sp_inst_18.INIT_RAM_12 = 256'h28BF57FD0015288028BF4C0028800010029E1C0000406802028102BF28000010;
defparam sp_inst_18.INIT_RAM_13 = 256'h028028BF29BF028028BF57FC00150067288028BF500229BF028028BF29BF0280;
defparam sp_inst_18.INIT_RAM_14 = 256'h500229BF028028BF29BF028028BF57FD001528BF02800015288028BF500229BF;
defparam sp_inst_18.INIT_RAM_15 = 256'h288028BF500129BF028028BF29BF028028BF57FD001528BF02800280288028BF;
defparam sp_inst_18.INIT_RAM_16 = 256'h02800015288028BF500129BF028028BF29BF028028BF57FD001528BF02800015;
defparam sp_inst_18.INIT_RAM_17 = 256'h001528BF02800015288028BF500129BF028028BF29BF028028BF57FC001528BF;
defparam sp_inst_18.INIT_RAM_18 = 256'h028028BF500129BF028028BF57FB0280500129BF028028BF29BF028028BF57FC;
defparam sp_inst_18.INIT_RAM_19 = 256'h028028BF29BF001002BF2800001028BF028028BF001C028028BF500029BF29BF;
defparam sp_inst_18.INIT_RAM_1A = 256'h53FD67FF02802800001028BF028028BF67FD02802800001028BF028028BF29BF;
defparam sp_inst_18.INIT_RAM_1B = 256'h29BF028028BF29BF001002BF2800001028BF028028BF001C028028BF500029BF;
defparam sp_inst_18.INIT_RAM_1C = 256'h028053FD67FF02802800001028BF028028BF67FD02802800001028BF028028BF;
defparam sp_inst_18.INIT_RAM_1D = 256'h0020028028BF400028BF57FA00152A3F57FA02805C000280283F5000034057FA;
defparam sp_inst_18.INIT_RAM_1E = 256'h28BF47FF29BF02BF28BF0340034003400340500029BF03AC14004400002A5C00;
defparam sp_inst_18.INIT_RAM_1F = 256'h0280298002BF4C000281288028800015001547FC2800001028BF28BF29BF0280;
defparam sp_inst_18.INIT_RAM_20 = 256'h028028800340040203800280298002BF4C0002802880001528BF29BF000029BF;
defparam sp_inst_18.INIT_RAM_21 = 256'h28BF29BF02802980298002BF4C00028028800340040203800280298002BF4C00;
defparam sp_inst_18.INIT_RAM_22 = 256'h02802980298002BF4C000280288028800340298028BF001557FF298028BF2980;
defparam sp_inst_18.INIT_RAM_23 = 256'h50000011288028BF288028BF6800288028BF288028BF298028BF001557FF29BF;
defparam sp_inst_18.INIT_RAM_24 = 256'h298002BF4C0002802880288000150010288028BF001128BF288028BF29BF02BF;
defparam sp_inst_18.INIT_RAM_25 = 256'h28BF29BF57FF001502BF500057FF001502BF57FE29BF29BF29BF29BF02802980;
defparam sp_inst_18.INIT_RAM_26 = 256'h0015004028BF29BF02802980298002BF4C00028028802880034057FE6BFF28BF;
defparam sp_inst_18.INIT_RAM_27 = 256'h0015001C03BD140028BF29BF02802980298002BF4C00028028802880034057FF;
defparam sp_inst_18.INIT_RAM_28 = 256'h57FF0015001C028F28BF29BF02802980298002BF4C00028028802880034057FF;
defparam sp_inst_18.INIT_RAM_29 = 256'h4400280029BF028028BF500029BF29BF0280298002BF4C000280288028800340;
defparam sp_inst_18.INIT_RAM_2A = 256'h28BF29BF02BF28BF00152A0028BF5BFF280029BF028028BF280028BF50000015;
defparam sp_inst_18.INIT_RAM_2B = 256'h29BF28800380157F29BF29BF29BF0280298002BF4C0002802880001500112A00;
defparam sp_inst_18.INIT_RAM_2C = 256'h006703400067004428BF290028BF006703410067004428BF29BF28800380157F;
defparam sp_inst_18.INIT_RAM_2D = 256'h28BF290028BF006703400067004428BF290028BF00670340006728BF290028BF;
defparam sp_inst_18.INIT_RAM_2E = 256'h028028800340290028BF006703400067004428BF290028BF0067034000670044;
defparam sp_inst_18.INIT_RAM_2F = 256'h28BF2900028028BF44002A0028BF680002802A0028BF29BF0280298002BF4C00;
defparam sp_inst_18.INIT_RAM_30 = 256'h002102802A0028BF29801410157F2900028028BF44002A0028BF680002802A00;
defparam sp_inst_18.INIT_RAM_31 = 256'h02802A0028BF001500400067002A5C00002102802A0028BF00400067002A5C00;
defparam sp_inst_18.INIT_RAM_32 = 256'h0380157F00150067002A5C00002102812A0028BF001500400067002A5C000021;
defparam sp_inst_18.INIT_RAM_33 = 256'h03402A0028BF001500400067002A5C00002102802A0028BF00402A0028BF2980;
defparam sp_inst_18.INIT_RAM_34 = 256'h02802980298002BF4C00028028800340298015000380157F29800380157F0015;
defparam sp_inst_18.INIT_RAM_35 = 256'h02BF4C00028028802880034057FE28BF500057FD28BF40002A3F293F29BF0015;
defparam sp_inst_18.INIT_RAM_36 = 256'h001728BF02802881157F440028BF29BF28BF6000028028BF29BF29BF02802980;
defparam sp_inst_18.INIT_RAM_37 = 256'h500029810015157F0015001728BF02802881157F500029810014157F00150014;
defparam sp_inst_18.INIT_RAM_38 = 256'h500029810014157F00150014001728BF02802881157F440028BF29BF02BF28BF;
defparam sp_inst_18.INIT_RAM_39 = 256'h0280298002BF4C0002802880034029810015157F0015001728BF02802881157F;
defparam sp_inst_18.INIT_RAM_3A = 256'h00150014001728BF02802881157F440028BF29BF28BF6000028028BF29BF29BF;
defparam sp_inst_18.INIT_RAM_3B = 256'h02BF28BF500029810015157F0015001728BF02802881157F500029810014157F;
defparam sp_inst_18.INIT_RAM_3C = 256'h2881157F500029810014157F00150014001728BF02802881157F440028BF29BF;
defparam sp_inst_18.INIT_RAM_3D = 256'h2A00157F0280298002BF4C0002802880034029810015157F0015001728BF0280;
defparam sp_inst_18.INIT_RAM_3E = 256'h28BF29BF29BF29BF0280298002BF4C00028028800340290000670380157F0067;
defparam sp_inst_18.INIT_RAM_3F = 256'h0380157F28800380157F2980001403BF15FB0380157F28800380157F40012880;

SP sp_inst_19 (
    .DO({sp_inst_19_dout_w[15:0],sp_inst_19_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_3}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_19.READ_MODE = 1'b0;
defparam sp_inst_19.WRITE_MODE = 2'b01;
defparam sp_inst_19.BIT_WIDTH = 16;
defparam sp_inst_19.BLK_SEL = 3'b001;
defparam sp_inst_19.RESET_MODE = "SYNC";
defparam sp_inst_19.INIT_RAM_00 = 256'h28BF5000298028BF00140014288028BF288028BF4400288028BF298000151404;
defparam sp_inst_19.INIT_RAM_01 = 256'h28BF288028BF298028BF0015288028BF288028BF298028BF0015288028BF2880;
defparam sp_inst_19.INIT_RAM_02 = 256'h298028BF0015288028BF288028BF5C000280288028BF298028BF001400142880;
defparam sp_inst_19.INIT_RAM_03 = 256'h298028BF0015288028BF288028BF298028BF00140014288028BF288028BF5000;
defparam sp_inst_19.INIT_RAM_04 = 256'h0280298002BF4C00028028800340298028BF00140014288028BF288028BF5000;
defparam sp_inst_19.INIT_RAM_05 = 256'h02BF4C00028028800340298028BF2980028028BF2980028028BF298028BF29BF;
defparam sp_inst_19.INIT_RAM_06 = 256'h298002BF4C00028028800340298028BF001528BF288028BF29BF29BF02802980;
defparam sp_inst_19.INIT_RAM_07 = 256'h0280288003402980001528BF157F0040001428BF29800396154A157F29BF0280;
defparam sp_inst_19.INIT_RAM_08 = 256'h02802980298002BF4C0002802880034029800396154A157F0280298002BF4C00;
defparam sp_inst_19.INIT_RAM_09 = 256'h29BF002A5C00002128BF288028BF2900028028BF29BF0388140029BF29BF29BF;
defparam sp_inst_19.INIT_RAM_0A = 256'h28BF2A0028BF290028BF0067004428BF290028BF006728BF29BF02BF004428BF;
defparam sp_inst_19.INIT_RAM_0B = 256'h28BF40002A0028BF290028BF0067001502BE006700152A0028BF006700152A00;
defparam sp_inst_19.INIT_RAM_0C = 256'h0280298002BF4C0002802880288003405402157F290028BF2A0028BF29000280;
defparam sp_inst_19.INIT_RAM_0D = 256'h290028BF2900028028BF2900028028BF2900028028BF2980039A140028BF29BF;
defparam sp_inst_19.INIT_RAM_0E = 256'h0067038100672A0028BF400028BF29BF29BF0280298002BF4C00028028800340;
defparam sp_inst_19.INIT_RAM_0F = 256'h02BF4C00028028800340290028BF0067001402BE00672A0028BF5000290028BF;
defparam sp_inst_19.INIT_RAM_10 = 256'h2880034029000280157F29002A3F28BF540128BF293F001529BF028029802980;
defparam sp_inst_19.INIT_RAM_11 = 256'h006728BF006728BF540128BF29BF29BF29BF02802980298002BF4C0002802880;
defparam sp_inst_19.INIT_RAM_12 = 256'h29BF02802980298002BF4C000280288028800340290028BF0067038000670015;
defparam sp_inst_19.INIT_RAM_13 = 256'h02A21C0000152A3F293F03802A3F40002A3F540028BF293F0015293F00150015;
defparam sp_inst_19.INIT_RAM_14 = 256'h02BE157F29002A3F28BF57E602A11C0000152A3F293F001402BF2A3F500057E6;
defparam sp_inst_19.INIT_RAM_15 = 256'h2A0028BF5000293F2A0028BF29BF0280298002BF4C0002802880288003402900;
defparam sp_inst_19.INIT_RAM_16 = 256'h2A3F293F2A0028BF29BF0280298002BF4C0002802880034047FF03402A3F293F;
defparam sp_inst_19.INIT_RAM_17 = 256'h2980298002BF4C00028028800340290028BF0067038000672A0028BF40000340;
defparam sp_inst_19.INIT_RAM_18 = 256'h2A3F293F02BE0067006F00442A7F297F035F2A7F293F0015297F001500150280;
defparam sp_inst_19.INIT_RAM_19 = 256'h00672A00157F57FE157F57FE157F001500152A3F57E5029D1C00001500152A3F;
defparam sp_inst_19.INIT_RAM_1A = 256'h001500672A7F57E5029D1C0000152A7F297F03432A7F57E5029D1C0064000000;
defparam sp_inst_19.INIT_RAM_1B = 256'h57FD157F00152A3F57E4029B1C006400000000672A00157F57FE157F57FD157F;
defparam sp_inst_19.INIT_RAM_1C = 256'h034057FE157F57FC157F028057E4029A1C006400000000672A00157F57FE157F;
defparam sp_inst_19.INIT_RAM_1D = 256'h006F00442A7F297F035F2A7F297F001502802980298002BF4C00028028802880;
defparam sp_inst_19.INIT_RAM_1E = 256'h157F57FD157F57FC157F001500152A3F57E402991C0000152A3F293F02BE0067;
defparam sp_inst_19.INIT_RAM_1F = 256'h2A7F297F03432A7F57E302981C0000152A7F57E302991C006400000000672A00;
defparam sp_inst_19.INIT_RAM_20 = 256'h02802A3F57E302971C006400000000672A00157F57FD157F57FB157F00150067;
defparam sp_inst_19.INIT_RAM_21 = 256'h157F0280028157E302961C006400000000672A00157F57FD157F57FC157F0015;
defparam sp_inst_19.INIT_RAM_22 = 256'h157F0280298002BF4C0002802880288000152A3F293F2A00157F57FC157F57FB;
defparam sp_inst_19.INIT_RAM_23 = 256'h03405FFF028028BF29BF28800380157F500029BF28800380157F298015000380;
defparam sp_inst_19.INIT_RAM_24 = 256'h0380157F500029BF28800380157F29BF29BF29BF0280298002BF4C0002802880;
defparam sp_inst_19.INIT_RAM_25 = 256'h28BF298028BF0380157F2980001403BF143F28BF157F5FFF028028BF29BF2880;
defparam sp_inst_19.INIT_RAM_26 = 256'h02BF4C00028028800340298002800380157F5000298002800380157F5C000280;
defparam sp_inst_19.INIT_RAM_27 = 256'h001403BF140000402A0028BF001500402A0028BF00402A0028BF29BF02802980;
defparam sp_inst_19.INIT_RAM_28 = 256'h034029800380157F001503402A0028BF0015001403BC140000402A0028BF0015;
defparam sp_inst_19.INIT_RAM_29 = 256'h00150014140100402A0028BF00402A0028BF29BF0280298002BF4C0002802880;
defparam sp_inst_19.INIT_RAM_2A = 256'h0380157F00152A0028BF0015037C00402A0028BF00150014140000402A0028BF;
defparam sp_inst_19.INIT_RAM_2B = 256'h140000402A0028BF00402A4028BF29BF0280298002BF4C000280288003402980;
defparam sp_inst_19.INIT_RAM_2C = 256'h2A0028BF0015036000402A0028BF00150014140000402A0028BF0015001403BF;
defparam sp_inst_19.INIT_RAM_2D = 256'h03402A0028BF0015034000402A0028BF0015034300402A0028BF0015034C0040;
defparam sp_inst_19.INIT_RAM_2E = 256'h28800380157F400028BF29BF0280298002BF4C000280288003402980157F0015;
defparam sp_inst_19.INIT_RAM_2F = 256'h0280288003402980001402B70380157F28800380157F5000298003880380157F;
defparam sp_inst_19.INIT_RAM_30 = 256'h006F037F006F288000100381157F001500402A7F297F00150280298002BF4C00;
defparam sp_inst_19.INIT_RAM_31 = 256'h288000100382157F001500402A7F297F00150280298002BF4C00028028800015;
defparam sp_inst_19.INIT_RAM_32 = 256'h034029800380157F2880157F0280298002BF4C00028028800015006F037F006F;
defparam sp_inst_19.INIT_RAM_33 = 256'h02BF4C0002802880034029800380157F2880157F0280298002BF4C0002802880;
defparam sp_inst_19.INIT_RAM_34 = 256'h2A3F037F288000100381157F001500402A3F293F0015293F0015001502802980;
defparam sp_inst_19.INIT_RAM_35 = 256'h298002BF4C000280288003402980001500100381157F001500402A3F00150040;
defparam sp_inst_19.INIT_RAM_36 = 256'h288000100382157F001500402A3F001500402A3F293F0015293F001500150280;
defparam sp_inst_19.INIT_RAM_37 = 256'h2980298002BF4C000280288003402980001500100381157F001500402A3F037F;
defparam sp_inst_19.INIT_RAM_38 = 256'h02802A7F297F02802A7F57FF001500152A3F00672A7F5000297F293F00150280;
defparam sp_inst_19.INIT_RAM_39 = 256'h293F0280293F0281293F001502812980298002BF4C0002802880288003406FFF;
defparam sp_inst_19.INIT_RAM_3A = 256'h293F0280293F0280293F293F028057FB001502BF293F0280293F0280293F0280;
defparam sp_inst_19.INIT_RAM_3B = 256'h293F0280293F0280293F293F0280293F0280297F03BF57FB001502BF293F02BF;
defparam sp_inst_19.INIT_RAM_3C = 256'h57FC028057FE00152A3F47FF03402880157F034057FD57FB001502BF293F293F;
defparam sp_inst_19.INIT_RAM_3D = 256'h001557FC0015006F28BF500029BF02812981298102BE4C000281288028800340;
defparam sp_inst_19.INIT_RAM_3E = 256'h29BF57DC02BC1C0067FF028028BF29BF028028BF29BF001002BF004028BF0015;
defparam sp_inst_19.INIT_RAM_3F = 256'h67FF028028BF29BF028028BF57DB02BA1C00001528BF001002BF004028BF5000;

SP sp_inst_20 (
    .DO({sp_inst_20_dout_w[15:0],sp_inst_20_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_4}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_20.READ_MODE = 1'b0;
defparam sp_inst_20.WRITE_MODE = 2'b01;
defparam sp_inst_20.BIT_WIDTH = 16;
defparam sp_inst_20.BLK_SEL = 3'b001;
defparam sp_inst_20.RESET_MODE = "SYNC";
defparam sp_inst_20.INIT_RAM_00 = 256'h4C00028128812881034057DB02BA1C0000152A3F293F0340006728800380157F;
defparam sp_inst_20.INIT_RAM_01 = 256'h0380157F2980288028BF0380157F29800380157F2980157F29BF0280298002BF;
defparam sp_inst_20.INIT_RAM_02 = 256'h00672A00157F4000288028BF29800015157F288028BF2880157F2980288028BF;
defparam sp_inst_20.INIT_RAM_03 = 256'h157F288028BF2880157F29800015157F288028BF2880157F290000670380157F;
defparam sp_inst_20.INIT_RAM_04 = 256'h028028BF29800388140028BF29BF0280298002BF4C0002802880034029800015;
defparam sp_inst_20.INIT_RAM_05 = 256'h28BF298003A2140028BF298003BC140028BF2980028028BF2980028028BF2980;
defparam sp_inst_20.INIT_RAM_06 = 256'h29800380157F2880157F400028BF29BF0280298002BF4C000280288003402980;
defparam sp_inst_20.INIT_RAM_07 = 256'h400028BF29BF0280298002BF4C0002802880034029800343157F2880157F5000;
defparam sp_inst_20.INIT_RAM_08 = 256'h157F2880157F5000290000670380157F00672A00157F29800380157F2880157F;
defparam sp_inst_20.INIT_RAM_09 = 256'h298002BF4C0002802880034029000067001402BF157F00672A00157F29800343;
defparam sp_inst_20.INIT_RAM_0A = 256'h02802880001528BF29BF500029BF02804000001428BF2880157F29BF29BF0280;
defparam sp_inst_20.INIT_RAM_0B = 256'h157F00672A000380157F2980001528BF157F2880157F29BF0280298002BF4C00;
defparam sp_inst_20.INIT_RAM_0C = 256'h28800015034029BF29BF0280298002BF4C000280288003402900006703800380;
defparam sp_inst_20.INIT_RAM_0D = 256'h1C0050015800028028BF5800028028BF29BF29BF02802980298002BF4C000280;
defparam sp_inst_20.INIT_RAM_0E = 256'h02811C000015001528800010004028BF02B91C00028028BF500029BF57D80281;
defparam sp_inst_20.INIT_RAM_0F = 256'h47FF001557E602B81C00001528800010004028BF02B91C0029BF028028BF57D8;
defparam sp_inst_20.INIT_RAM_10 = 256'h001557E628BF001528800010004028BF02B71C00500029BF29BF288028BF5001;
defparam sp_inst_20.INIT_RAM_11 = 256'h28BF02B61C0028800010004028BF02B61C0028800010004028BF02B71C004400;
defparam sp_inst_20.INIT_RAM_12 = 256'h28BF02B51C0029BF028028BF500057D702BD1C00001500150015288000100040;
defparam sp_inst_20.INIT_RAM_13 = 256'h001528800010004028BF02B41C0047FF001557E502B41C000015288000100040;
defparam sp_inst_20.INIT_RAM_14 = 256'h001500150340500057D602BC1C00500057D602BC1C004400001557E502B41C00;
defparam sp_inst_20.INIT_RAM_15 = 256'h29BF03BF1400298002800380157F57DB02812980298002BF4C00028028802880;
defparam sp_inst_20.INIT_RAM_16 = 256'h500029BF03AC140057DE02BA1C0047FF29BF02BF28BF03400340034003405000;
defparam sp_inst_20.INIT_RAM_17 = 256'h140057DE02B91C0028BF29BF02B91C0047FF29BF02BF28BF0340034003400340;
defparam sp_inst_20.INIT_RAM_18 = 256'h1C00028029BF0389148847FF29BF02BF28BF0340034003400340500029BF03AC;
defparam sp_inst_20.INIT_RAM_19 = 256'h29BF028047FF29BF02BF28BF0340034003400340500029BF03AC140057DD02B8;
defparam sp_inst_20.INIT_RAM_1A = 256'h29BF02BF28BF0340034003400340500029BF03AC140057DD02B71C00001528BF;
defparam sp_inst_20.INIT_RAM_1B = 256'h0340034003400340500029BF03BF140057E857E60280028057E60280028047FF;
defparam sp_inst_20.INIT_RAM_1C = 256'h28BF0340034003400340500029BF03BF140057E70280028047FF29BF02BF28BF;
defparam sp_inst_20.INIT_RAM_1D = 256'h02BF4C0002802880001500150280298002BF53FF57E70280001547FF29BF02BF;
defparam sp_inst_20.INIT_RAM_1E = 256'h5000028057D402B31C006400028028BF6400028028BF29BF29BF028029802980;
defparam sp_inst_20.INIT_RAM_1F = 256'h00152880028028BF500029BF02805C00028028BF29BF540200152880028028BF;
defparam sp_inst_20.INIT_RAM_20 = 256'h28BF57D302B11C000015001028BF28BF4400034028BF500029BF29BF00155402;
defparam sp_inst_20.INIT_RAM_21 = 256'h0015001563FF28BF28BF29BF028028BF57D302B11C00001500672A00001028BF;
defparam sp_inst_20.INIT_RAM_22 = 256'h6400028028BF6400028028BF29BF29BF02802980298002BF4C00028028802880;
defparam sp_inst_20.INIT_RAM_23 = 256'h29BF02805C00028028BF29BF540100152880028028BF5000028057D302AF1C00;
defparam sp_inst_20.INIT_RAM_24 = 256'h0015004028BF4400034028BF500029BF29BF0015540100152880028028BF5000;
defparam sp_inst_20.INIT_RAM_25 = 256'h57D202AD1C0000152880001028BF0015004028BF57D202AE1C000015001028BF;
defparam sp_inst_20.INIT_RAM_26 = 256'h02802980298002BF4C000280288028800015001563FF28BF28BF29BF028028BF;
defparam sp_inst_20.INIT_RAM_27 = 256'h29BF540000152880028028BF5000028057D102AC1C005800028028BF29BF29BF;
defparam sp_inst_20.INIT_RAM_28 = 256'h4C000280288028800015001529002A3F28BF293F0015540000152880028028BF;
defparam sp_inst_20.INIT_RAM_29 = 256'h028028BF5000028057D102AA1C005800028028BF29BF29BF02802980298002BF;
defparam sp_inst_20.INIT_RAM_2A = 256'h288000150015298028BF28BF29BF540000152880028028BF29BF540000152880;
defparam sp_inst_20.INIT_RAM_2B = 256'h2A00028028BF5C0002802A0028BF29BF29BF02802980298002BF4C0002802880;
defparam sp_inst_20.INIT_RAM_2C = 256'h5C0002802A0028BF500029BF028029BF02805C0002812A00028028BF58000281;
defparam sp_inst_20.INIT_RAM_2D = 256'h028028BF29BF2A00001028BF28BF500129BF028029BF500129BF028029BF0280;
defparam sp_inst_20.INIT_RAM_2E = 256'h28BF28BF6800028028BF6C00028028BF50015800028028BF5800028028BF5800;
defparam sp_inst_20.INIT_RAM_2F = 256'h28BF001C28BF28BF6800028128BF6C00028128BF500029BF02BF001028BF001C;
defparam sp_inst_20.INIT_RAM_30 = 256'h02BF001028BF001C28BF28BF6800028128BF6C00028128BF500029BF02BE0010;
defparam sp_inst_20.INIT_RAM_31 = 256'h28BF28BF6C0028BF028028BF6C00028028BF5000500057CF02A31C00500029BF;
defparam sp_inst_20.INIT_RAM_32 = 256'h001028BF28BF29BF028028BF034057CF02A21C00500029BF02BF001028BF001C;
defparam sp_inst_20.INIT_RAM_33 = 256'h028028BF29BF29BF02802980298002BF4C00028028802880001528BF47FE2A00;
defparam sp_inst_20.INIT_RAM_34 = 256'h00152880028028BF29BF57FD00152880028028BF5000028057CE02A11C005800;
defparam sp_inst_20.INIT_RAM_35 = 256'h28800015001557CE02A01C0057EB28BF28BF028057CE02A01C0057EB29BF57FD;
defparam sp_inst_20.INIT_RAM_36 = 256'h57CE029F1C0000152880157F57CE02A01C0002802980298002BF4C0002802880;
defparam sp_inst_20.INIT_RAM_37 = 256'h029F1C0057CD029F1C00001528800380157F57CD029F1C00001528800380157F;
defparam sp_inst_20.INIT_RAM_38 = 256'h00100382157F0015004028BF288000100381157F0015004028BF500029BF57CD;
defparam sp_inst_20.INIT_RAM_39 = 256'h28800015001567FF028028BF29BF028028BF57CD029E1C0028BF001500152880;
defparam sp_inst_20.INIT_RAM_3A = 256'h28BF500029BF57CD029F1C0057CD029E1C0002802980298002BF4C0002802880;
defparam sp_inst_20.INIT_RAM_3B = 256'h029E1C0067FF028028BF29BF028028BF57CC029E1C000015001557ED0015006F;
defparam sp_inst_20.INIT_RAM_3C = 256'h28BF29BF028028BF57CC029D1C000015001557ED0015006F28BF500029BF57CC;
defparam sp_inst_20.INIT_RAM_3D = 256'h028028BF29BF29BF02802980298002BF4C000280288028800015001567FF0280;
defparam sp_inst_20.INIT_RAM_3E = 256'h1C005002028057CC029B1C005800028028BF4400001557DA029B1C0000152880;
defparam sp_inst_20.INIT_RAM_3F = 256'h2880028028BF500257EE00152A3F293F001557FA00152880028028BF57CC029B;

SP sp_inst_21 (
    .DO({sp_inst_21_dout_w[15:0],sp_inst_21_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_5}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_21.READ_MODE = 1'b0;
defparam sp_inst_21.WRITE_MODE = 2'b01;
defparam sp_inst_21.BIT_WIDTH = 16;
defparam sp_inst_21.BLK_SEL = 3'b001;
defparam sp_inst_21.RESET_MODE = "SYNC";
defparam sp_inst_21.INIT_RAM_00 = 256'h029A1C004000006700140067024003C028BF00670240001557DA029A1C000015;
defparam sp_inst_21.INIT_RAM_01 = 256'h57CB02991C004400001557D902991C0000152880028028BF500157EF57EC57CB;
defparam sp_inst_21.INIT_RAM_02 = 256'h001500152A3F2A3F5000293F5C00028028BF293F001557FA00152880028028BF;
defparam sp_inst_21.INIT_RAM_03 = 256'h57F900152880028028BF5C00028028BF50016FFF02802A3F293F02802A3F57EC;
defparam sp_inst_21.INIT_RAM_04 = 256'h2880028028BF5000028057CA02971C00500057EB001500152A3F2A3F293F0015;
defparam sp_inst_21.INIT_RAM_05 = 256'h02961C004000006700140067024003C028BF00670240001557D902971C000015;
defparam sp_inst_21.INIT_RAM_06 = 256'h024003C028BF00670240001557D802961C0000152880028028BF500057EB57CA;
defparam sp_inst_21.INIT_RAM_07 = 256'h00155000028057C902951C0057C902951C00500057FC57FB4000006700140067;
defparam sp_inst_21.INIT_RAM_08 = 256'h028028BE57C902961C0029BE29BE02812981298102BE4C000280288028800015;
defparam sp_inst_21.INIT_RAM_09 = 256'h29BF57F800152880028028BE5000028057C902961C0057EF001557EF00156000;
defparam sp_inst_21.INIT_RAM_0A = 256'h28BF57EE001502BF29BF57F800152880028028BE29BF57F800152880028028BE;
defparam sp_inst_21.INIT_RAM_0B = 256'h001557ED001502BF29BF001C0388140028BF29BF001C03BC140028BF29BF0040;
defparam sp_inst_21.INIT_RAM_0C = 256'h28BF57C802931C0028BF29BF29BF02802980298002BF4C000281288128810015;
defparam sp_inst_21.INIT_RAM_0D = 256'h140128BF29BF57F700152880028028BF5000028057C802931C0057CD60000280;
defparam sp_inst_21.INIT_RAM_0E = 256'h29BF29BF02802980298002BF4C000280288028800015001557CD0015001C038F;
defparam sp_inst_21.INIT_RAM_0F = 256'h028028BF29BF57F600152880028028BF5000028057C702911C006000028028BF;
defparam sp_inst_21.INIT_RAM_10 = 256'h028028BF500057C702911C0028BF57D528BF5C00028028BF29BF57F600152880;
defparam sp_inst_21.INIT_RAM_11 = 256'h02901C0028BF57D528BF5C00028028BF500057C702901C0028BF57D528BF5C00;
defparam sp_inst_21.INIT_RAM_12 = 256'h29BF02802980298002BF4C000280288028800015001557C7028E1C00500057C7;
defparam sp_inst_21.INIT_RAM_13 = 256'h5000028057C6028F1C0057CC00156000028028BF57CB57C6028F1C0028BF29BF;
defparam sp_inst_21.INIT_RAM_14 = 256'h02BF4C000280288028800015001557BC57CC28BF29BF57F500152880028028BF;
defparam sp_inst_21.INIT_RAM_15 = 256'h500002BF57C6028D1C006C0002802A3F6C0002802A3F293F0015028029802980;
defparam sp_inst_21.INIT_RAM_16 = 256'h028C1C0029BD29BD028229822982298202BD4C00028028802880001503402A3F;
defparam sp_inst_21.INIT_RAM_17 = 256'h001528BD2880028028BD29BE29BE29BD29BD288028802880288002911C0057C6;
defparam sp_inst_21.INIT_RAM_18 = 256'h57C5028C1C0057C5028C1C0057C5028B1C0057C5028B1C004400001557D40015;
defparam sp_inst_21.INIT_RAM_19 = 256'h028C1C005800028028BD4402001557D30015001528BD2880028028BD50060015;
defparam sp_inst_21.INIT_RAM_1A = 256'h001C0280001557FE00152A0028BF29BF288028BD29BF288028BD5006028057C5;
defparam sp_inst_21.INIT_RAM_1B = 256'h001C0280001557FE00152A00028028BF29BF0010001557FE00152A00028028BF;
defparam sp_inst_21.INIT_RAM_1C = 256'h001C0280001557FE00152A00028028BF29BF0010001557FE00152A00028028BF;
defparam sp_inst_21.INIT_RAM_1D = 256'h28BF001C0280001557FD00152A0028BF29BF0010001557FD00152A00028028BF;
defparam sp_inst_21.INIT_RAM_1E = 256'h28BF001C0280001557FD00152A00028028BF29BF0010001557FD00152A000280;
defparam sp_inst_21.INIT_RAM_1F = 256'h28BF001C0280001557FD00152A00028028BF29BF0010001557FD00152A000280;
defparam sp_inst_21.INIT_RAM_20 = 256'h28BF6800028028BF400028BF6800028028BF29BF0010001557FD00152A000280;
defparam sp_inst_21.INIT_RAM_21 = 256'h6C00028028BF6800028028BF6800028028BF6800028028BF5C00028028BF4000;
defparam sp_inst_21.INIT_RAM_22 = 256'h006728BF293D006728BF5003028057C302841C00400028BF29BF001550000280;
defparam sp_inst_21.INIT_RAM_23 = 256'h0015001502BD293D006728BF293D006728BF293D006728BF293D006728BF293D;
defparam sp_inst_21.INIT_RAM_24 = 256'h02811C005800028028BD4402001557D10015001528BE2880028028BD500357D4;
defparam sp_inst_21.INIT_RAM_25 = 256'h001C0280001557FB00152A0028BF29BF288028BD29BF288028BD5003028057C2;
defparam sp_inst_21.INIT_RAM_26 = 256'h001C0280001557FB00152A00028028BF29BF0010001557FB00152A00028028BF;
defparam sp_inst_21.INIT_RAM_27 = 256'h28BF001C0280001557FB00152A0028BF29BE0010001557FB00152A00028028BF;
defparam sp_inst_21.INIT_RAM_28 = 256'h28BF001C0280001557FB00152A00028028BF29BE0010001557FB00152A000280;
defparam sp_inst_21.INIT_RAM_29 = 256'h28BF001C0280001557FA00152A00028028BF29BE0010001557FA00152A000280;
defparam sp_inst_21.INIT_RAM_2A = 256'h28BE6800028028BE400028BF6800028028BF29BE0010001557FA00152A000280;
defparam sp_inst_21.INIT_RAM_2B = 256'h6C00028028BE6800028028BE6800028028BE6800028028BE5C00028028BF4000;
defparam sp_inst_21.INIT_RAM_2C = 256'h006728BE293D006728BE5001028057C002BA1C00400028BE29BE001550000280;
defparam sp_inst_21.INIT_RAM_2D = 256'h28BE2880028028BD50010015293D006728BF293D006728BE293D006728BE293D;
defparam sp_inst_21.INIT_RAM_2E = 256'h006700120394140028BE29BE57EF00152880028028BD4400001557CE00150015;
defparam sp_inst_21.INIT_RAM_2F = 256'h004428BE5000028057BF02B71C00400000670015006703C00012038D140028BE;
defparam sp_inst_21.INIT_RAM_30 = 256'h57D00280001502BD57BF02B61C005800028028BD5000001529BE034028BE29BE;
defparam sp_inst_21.INIT_RAM_31 = 256'h1C0028BE28BE28BE29BE2A3D29BE2A3D29BE2A3D29BE2A3D29BE2A3D29BE2A3D;
defparam sp_inst_21.INIT_RAM_32 = 256'h02BF4C0002822882288228820015001557BF02B51C0028BE28BE28BE57BF02B5;
defparam sp_inst_21.INIT_RAM_33 = 256'h57BE02B51C0057D56000028028BF57BE02B51C0028BF29BF29BF028029802980;
defparam sp_inst_21.INIT_RAM_34 = 256'h4C000280288028800015001557D428BF29BF57ED00152880028028BF50000280;
defparam sp_inst_21.INIT_RAM_35 = 256'h28800015034057D4157F001502BF57D5001502BF29BF29BF02802980298002BF;
defparam sp_inst_21.INIT_RAM_36 = 256'h028057BE02B21C005800028028BF29BF29BF02802980298002BF4C0002802880;
defparam sp_inst_21.INIT_RAM_37 = 256'h57EC00152880028028BF293F001557EC00152880028028BF57BE02AC1C005000;
defparam sp_inst_21.INIT_RAM_38 = 256'h0000001500002A3F000000402A3F293F001557EC00152880028028BF293F0015;
defparam sp_inst_21.INIT_RAM_39 = 256'h57D7001500152A7F2A3F57BD02B01C0000152A7F57BD02B11C0000152A3F297F;
defparam sp_inst_21.INIT_RAM_3A = 256'h1C005800028028BF29BF29BF02802980298002BF4C0002802880288000150015;
defparam sp_inst_21.INIT_RAM_3B = 256'h29BF57EB00152880028028BF29BF57EB00152880028028BF5000028057BD02AF;
defparam sp_inst_21.INIT_RAM_3C = 256'h00152A7F297F0015006F0343006F28BF006F001403BE1400006F0040006F28BF;
defparam sp_inst_21.INIT_RAM_3D = 256'h298002BF4C000280288028800015001557BC02AD1C0000152A3F293F001557D8;
defparam sp_inst_21.INIT_RAM_3E = 256'h29BF57EB00152880028028BF29BF57EB00152880028028BF29BF29BF02812980;
defparam sp_inst_21.INIT_RAM_3F = 256'h29BF0015500002806400028028BF6400028028BF6800028028BF6800028028BF;

SP sp_inst_22 (
    .DO({sp_inst_22_dout_w[15:0],sp_inst_22_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_6}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_22.READ_MODE = 1'b0;
defparam sp_inst_22.WRITE_MODE = 2'b01;
defparam sp_inst_22.BIT_WIDTH = 16;
defparam sp_inst_22.BLK_SEL = 3'b001;
defparam sp_inst_22.RESET_MODE = "SYNC";
defparam sp_inst_22.INIT_RAM_00 = 256'h1C0057BB02AB1C0057BB02AA1C00400028BF29BF001557EA00152880028028BF;
defparam sp_inst_22.INIT_RAM_01 = 256'h2980001028BF0381157F004028BF5000298014000380157F5000028057BB02AC;
defparam sp_inst_22.INIT_RAM_02 = 256'h00150044001C03B428BF29BF28800381157F298003840381157F28800381157F;
defparam sp_inst_22.INIT_RAM_03 = 256'h001403BF15FF0380157F28800380157F47FF28BF29BF02BF28BF57BB02AA1C00;
defparam sp_inst_22.INIT_RAM_04 = 256'h5800028028BF29BF29BF02802980298002BF4C00028128802880001500152980;
defparam sp_inst_22.INIT_RAM_05 = 256'h157F2880157F440028BF29BF57E900152880028028BF5001028057BA02A81C00;
defparam sp_inst_22.INIT_RAM_06 = 256'h157F50005800028028BF400028BF5800028028BF6800028028BF298000151400;
defparam sp_inst_22.INIT_RAM_07 = 256'h2880157F2980001403BF15F9157F2880157F50002980001403BF15F9157F2880;
defparam sp_inst_22.INIT_RAM_08 = 256'h1406157F2880157F2980001403BF15F9157F2880157F5000298000151404157F;
defparam sp_inst_22.INIT_RAM_09 = 256'h288000150015298003A00380157F5000028057B902A51C005000034029800015;
defparam sp_inst_22.INIT_RAM_0A = 256'h157F298002BF0380157F298002BF0380157F02802980298002BF4C0002802880;
defparam sp_inst_22.INIT_RAM_0B = 256'h1C0057CF298000151540157F001403BF140028BF500029BF157E298002800380;
defparam sp_inst_22.INIT_RAM_0C = 256'h28BF2980288028BF0015001015FE28BF500029BF28BF29801480157F57B802A3;
defparam sp_inst_22.INIT_RAM_0D = 256'h028228BF2980001515C0157F001403BF140028BF67FF28BF028128BF29BF0280;
defparam sp_inst_22.INIT_RAM_0E = 256'h2880001015FE28BF288028BF500029BF28BF500029BF157E6BFF157E28BF29BF;
defparam sp_inst_22.INIT_RAM_0F = 256'h157E28BF29BF028228BF67FF28BF028128BF29BF028028BF57B8029F1C005800;
defparam sp_inst_22.INIT_RAM_10 = 256'h5800028028BF29BF29BF02802980298002BF4C00028028802880001500156BFF;
defparam sp_inst_22.INIT_RAM_11 = 256'h57BA157F5C00028028BF29BF57E600152880028028BF5000028057B7029E1C00;
defparam sp_inst_22.INIT_RAM_12 = 256'h28802880001500155000028057B7029C1C00500057BA157F5C00028028BF5000;
defparam sp_inst_22.INIT_RAM_13 = 256'h001557B229000280157F29000281157F29BF29BF02802980298002BF4C000280;
defparam sp_inst_22.INIT_RAM_14 = 256'h02812980298002BF4C000280288028800015034057B6029B1C0000152A7F297F;
defparam sp_inst_22.INIT_RAM_15 = 256'h29BF57E500152880028028BF5000028057B6029A1C005800028028BF29BF29BF;
defparam sp_inst_22.INIT_RAM_16 = 256'h001028BF28BF500029BF29BF004028BF500029BF29BF028857B6029A1C0029BF;
defparam sp_inst_22.INIT_RAM_17 = 256'h1C006FFF028328BF29BF028028BF290000672A00001028BF28BF00150010157E;
defparam sp_inst_22.INIT_RAM_18 = 256'h1C006BFF28BF28BF29BF028028BF57B2001528BF0284001028BF28BF57B50298;
defparam sp_inst_22.INIT_RAM_19 = 256'h028028BF29BF29BF02812980298002BF4C000281288028800015001557B50297;
defparam sp_inst_22.INIT_RAM_1A = 256'h57B502961C0029BF29BF57E400152880028028BF5001028057B502961C005800;
defparam sp_inst_22.INIT_RAM_1B = 256'h500029BF57B2001528BF0284001028BF28BF29BF004028BF500029BF29BF0288;
defparam sp_inst_22.INIT_RAM_1C = 256'h2A00001028BF28BF580000672A000010157E001028BF28BF2A00001028BF28BF;
defparam sp_inst_22.INIT_RAM_1D = 256'h28BF29BF028028BF500057B402931C00001500150010157E001028BF28BF0015;
defparam sp_inst_22.INIT_RAM_1E = 256'h0015001557B402911C006BFF28BF28BF29BF028028BF57B402921C006FFF0283;
defparam sp_inst_22.INIT_RAM_1F = 256'h57B302911C005800028028BF29BF29BF02802980298002BF4C00028128802880;
defparam sp_inst_22.INIT_RAM_20 = 256'h0010140028BF57AF28BF57B302911C0029BF57E200152880028028BF50000280;
defparam sp_inst_22.INIT_RAM_21 = 256'h29BF29BF29BF29BF02812980298002BF4C000280288028800015001557AF0015;
defparam sp_inst_22.INIT_RAM_22 = 256'h57AF28BF57B3028C1C0000152A7F297F001557AE29000280157F29000281157F;
defparam sp_inst_22.INIT_RAM_23 = 256'h29BF29BF004028BF500029BF29BF028857B2028F1C0057AF00150010140028BF;
defparam sp_inst_22.INIT_RAM_24 = 256'h29BF028028BF290000672A00001028BF28BF00150010157E001028BF28BF5000;
defparam sp_inst_22.INIT_RAM_25 = 256'h29BF028028BF57B2028A1C0057AF001528BF0284001028BF28BF6FFF028328BF;
defparam sp_inst_22.INIT_RAM_26 = 256'h29BF004028BF500029BF29BF028857B2028C1C0057B2028C1C006BFF28BF28BF;
defparam sp_inst_22.INIT_RAM_27 = 256'h001028BF28BF2A00001028BF28BF500029BF57AF001528BF0284001028BF28BF;
defparam sp_inst_22.INIT_RAM_28 = 256'h00150010157E001028BF28BF00152A00001028BF28BF580000672A000010157E;
defparam sp_inst_22.INIT_RAM_29 = 256'h028028BF57B102861C006FFF028328BF29BF028028BF500057B102881C000015;
defparam sp_inst_22.INIT_RAM_2A = 256'h2980298002BF4C000281288028800015001557B102881C006BFF28BF28BF29BF;
defparam sp_inst_22.INIT_RAM_2B = 256'h0380140057C6001502BF57A80380157F0280001557A80380157F028000150280;
defparam sp_inst_22.INIT_RAM_2C = 256'h288028800015034057C40380157F001502BF29BF028029BF028029BF028029BF;
defparam sp_inst_22.INIT_RAM_2D = 256'h02BF4C000280288028800015001557FF29BF29BF02802980298002BF4C000280;
defparam sp_inst_22.INIT_RAM_2E = 256'h29BF29BF02802980298002BF4C00028028800015001529BF29BF29BF02802980;
defparam sp_inst_22.INIT_RAM_2F = 256'h29BF6BFF140028BF29BF028028BF29800010150028BF500029BF57B002841C00;
defparam sp_inst_22.INIT_RAM_30 = 256'h140028BF29BF028028BF2980288000150010150028BF00150010157C28BF5000;
defparam sp_inst_22.INIT_RAM_31 = 256'h28800010150028BF580028800010157C28BF28800010150028BF500029BF6BFF;
defparam sp_inst_22.INIT_RAM_32 = 256'h6BFF140028BF29BF028028BF57AF02811C0028BF0015001528800010157C28BF;
defparam sp_inst_22.INIT_RAM_33 = 256'h1C00028002861C0002802980298002BF4C00028028802880001500154C001500;
defparam sp_inst_22.INIT_RAM_34 = 256'h1C0002802980298002BF4C00028028802880034057C40380157F028057AE0280;
defparam sp_inst_22.INIT_RAM_35 = 256'h298002BF4C00028028802880034057C40380157F028057AE02BF1C0002800285;
defparam sp_inst_22.INIT_RAM_36 = 256'h028028802880034057C30380157F028057AE02BD1C00028002851C0002802980;
defparam sp_inst_22.INIT_RAM_37 = 256'h034057C30380157F028057AD02BC1C00028002841C0002802980298002BF4C00;
defparam sp_inst_22.INIT_RAM_38 = 256'h157F028057AD02BB1C00028002831C0002802980298002BF4C00028028802880;
defparam sp_inst_22.INIT_RAM_39 = 256'h02BA1C00028002821C0002802980298002BF4C00028028802880034057C30380;
defparam sp_inst_22.INIT_RAM_3A = 256'h02811C0002802980298002BF4C00028028802880034057C20380157F028057AD;
defparam sp_inst_22.INIT_RAM_3B = 256'h2980298002BF4C00028028802880034057C20380157F028157AD02B91C000280;
defparam sp_inst_22.INIT_RAM_3C = 256'h4C00028028802880034057C20380157F028257AC02B71C00028002811C000280;
defparam sp_inst_22.INIT_RAM_3D = 256'h2880034057C20380157F028457AC02B61C00028102801C0002802980298002BF;
defparam sp_inst_22.INIT_RAM_3E = 256'h0380157F028857AC02B51C00028102BF1C0002802980298002BF4C0002802880;
defparam sp_inst_22.INIT_RAM_3F = 256'h57AB02B41C00028102BE1C0002802980298002BF4C00028028802880034057C1;

SP sp_inst_23 (
    .DO({sp_inst_23_dout_w[15:0],sp_inst_23_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_7}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_23.READ_MODE = 1'b0;
defparam sp_inst_23.WRITE_MODE = 2'b01;
defparam sp_inst_23.BIT_WIDTH = 16;
defparam sp_inst_23.BLK_SEL = 3'b001;
defparam sp_inst_23.RESET_MODE = "SYNC";
defparam sp_inst_23.INIT_RAM_00 = 256'h028102BD1C0002802980298002BF4C00028028802880034057C10380157F0290;
defparam sp_inst_23.INIT_RAM_01 = 256'h02802980298002BF4C00028028802880034057C10380157F03A057AB02B31C00;
defparam sp_inst_23.INIT_RAM_02 = 256'h02BF4C00028028802880034057C00380157F140057AB02B11C00028102BD1C00;
defparam sp_inst_23.INIT_RAM_03 = 256'h28802880034057C00380157F140057AA02B01C00028102BC1C00028029802980;
defparam sp_inst_23.INIT_RAM_04 = 256'h57C00380157F140057AA02AF1C00028102BB1C0002802980298002BF4C000280;
defparam sp_inst_23.INIT_RAM_05 = 256'h140057AA02AE1C00028102BA1C0002802980298002BF4C000280288028800340;
defparam sp_inst_23.INIT_RAM_06 = 256'h1C00028102B91C0002802980298002BF4C00028028802880034057BF0380157F;
defparam sp_inst_23.INIT_RAM_07 = 256'h1C0002802980298002BF4C00028028802880034057BF0380157F140057AA02AD;
defparam sp_inst_23.INIT_RAM_08 = 256'h298002BF4C00028028802880034057BF0380157F140057A902AC1C00028102B8;
defparam sp_inst_23.INIT_RAM_09 = 256'h028028802880034057BF0380157F140057A902AA1C00028102B81C0002802980;
defparam sp_inst_23.INIT_RAM_0A = 256'h034057BE0380157F140057A902A91C00028202B71C0002802980298002BF4C00;
defparam sp_inst_23.INIT_RAM_0B = 256'h157F140057A802A81C00028202B61C0002802980298002BF4C00028028802880;
defparam sp_inst_23.INIT_RAM_0C = 256'h02A71C00028202B51C0002802980298002BF4C00028028802880034057BE0380;
defparam sp_inst_23.INIT_RAM_0D = 256'h02B41C0002802980298002BF4C00028028802880034057BE0380157F140057A8;
defparam sp_inst_23.INIT_RAM_0E = 256'h2980298002BF4C00028028802880034057BD0380157F140057A802A61C000282;
defparam sp_inst_23.INIT_RAM_0F = 256'h4C00028028802880034057BD0380157F140157A702A41C00028202B41C000280;
defparam sp_inst_23.INIT_RAM_10 = 256'h2880034057BD0380157F140257A702A31C00028202B31C0002802980298002BF;
defparam sp_inst_23.INIT_RAM_11 = 256'h0380157F140457A702A21C00028202B21C0002802980298002BF4C0002802880;
defparam sp_inst_23.INIT_RAM_12 = 256'h57A702A11C00028202B11C0002802980298002BF4C00028028802880034057BC;
defparam sp_inst_23.INIT_RAM_13 = 256'h028202B01C0002802980298002BF4C00028028802880034057BC0380157F1408;
defparam sp_inst_23.INIT_RAM_14 = 256'h02802980298002BF4C00028028802880034057BC0380157F141057A602A01C00;
defparam sp_inst_23.INIT_RAM_15 = 256'h02BF4C00028028802880034057BC0380157F142057A6029E1C00028202B01C00;
defparam sp_inst_23.INIT_RAM_16 = 256'h28802880034057BB0380157F144057A6029D1C00028202AF1C00028029802980;
defparam sp_inst_23.INIT_RAM_17 = 256'h57BB0380157F148057A5029C1C00028302AE1C0002802980298002BF4C000280;
defparam sp_inst_23.INIT_RAM_18 = 256'h150057A5029B1C00028302AD1C0002802980298002BF4C000280288028800340;
defparam sp_inst_23.INIT_RAM_19 = 256'h298014020380157F02802980298002BF4C00028028802880034057BB0380157F;
defparam sp_inst_23.INIT_RAM_1A = 256'h28BF28BF29BF28800380157F29BF28800380157F57A502991C00028302AC1C00;
defparam sp_inst_23.INIT_RAM_1B = 256'h28800010004028BF029B1C0040000340001728BF28BF500029BF034029BF0014;
defparam sp_inst_23.INIT_RAM_1C = 256'h02802980298002BF4C0002802880288003406FFF028028BF29BF028028BF4C00;
defparam sp_inst_23.INIT_RAM_1D = 256'h298002BF4C00028028802880034057BA29BF28800380157F298014000380157F;
defparam sp_inst_23.INIT_RAM_1E = 256'h157F293F0340006728800380157F297F037F006F004428800380157F02802980;
defparam sp_inst_23.INIT_RAM_1F = 256'h028028802880034057A302951C0000152A7F298002800380157F298014000380;
defparam sp_inst_23.INIT_RAM_20 = 256'h4C00028028800340293F2A000380157F298014000380157F0280298002BF4C00;
defparam sp_inst_23.INIT_RAM_21 = 256'h14010380157F28800380157F29BF0340004428800380157F02802980298002BF;
defparam sp_inst_23.INIT_RAM_22 = 256'h157F57A302931C004C002880001002971C00004028BF6800028028BF29800014;
defparam sp_inst_23.INIT_RAM_23 = 256'h50002980001403BF15FF0380157F28800380157F57A202931C00500029800380;
defparam sp_inst_23.INIT_RAM_24 = 256'h03402A3F293F2A000380157F02802980298002BF4C0002802880288003400340;
defparam sp_inst_23.INIT_RAM_25 = 256'h029A1CC72980029A1CC70015006702402880029A1CC74000001557C902844000;
defparam sp_inst_23.INIT_RAM_26 = 256'h157F5000293F28800380157F29BF400003402A3F57C9028457B4028000152880;
defparam sp_inst_23.INIT_RAM_27 = 256'h0280157F29BF400028BF500029BF028029800280157F5C00028028BF29BF2880;
defparam sp_inst_23.INIT_RAM_28 = 256'h157F400003402A3F43FF0340283F293F28800380157F298028BF157F50002980;
defparam sp_inst_23.INIT_RAM_29 = 256'h02802980298002BF4C000280288028800340290002BF0380157F290002800380;
defparam sp_inst_23.INIT_RAM_2A = 256'h0000000000000000000000004C00028028802880034057A657A1028C1C0057A6;
defparam sp_inst_23.INIT_RAM_2B = 256'h1C001C001C001C001C001C001C001C001C00000065646139363532310A21656B;
defparam sp_inst_23.INIT_RAM_2C = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_23.INIT_RAM_2D = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_23.INIT_RAM_2E = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_23.INIT_RAM_2F = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_23.INIT_RAM_30 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_23.INIT_RAM_31 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_23.INIT_RAM_32 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_23.INIT_RAM_33 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_23.INIT_RAM_34 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_23.INIT_RAM_35 = 256'h72201C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_23.INIT_RAM_36 = 256'h303D6441636944200000783278306464736E742000000A0D3025207261206965;
defparam sp_inst_23.INIT_RAM_37 = 256'h2064722000007830646400002D2D2D6B206F2D2D000078323020617454207832;
defparam sp_inst_23.INIT_RAM_38 = 256'h505500006F440000006400007830646400006B636F6E000032253D72415F6976;
defparam sp_inst_23.INIT_RAM_39 = 256'h093039303009093635303009093231303009000020746F4300006F44754D0000;
defparam sp_inst_23.INIT_RAM_3A = 256'h2D2D006C746E000064330000643200006C617553000064340000615661420000;
defparam sp_inst_23.INIT_RAM_3B = 256'h756400003E6D3C2064642031000000000000697800007469000025783A655479;
defparam sp_inst_23.INIT_RAM_3C = 256'h706C0064772065726120756400003E6D3C206464203400000065622065726120;
defparam sp_inst_23.INIT_RAM_3D = 256'h6F6D005D756C3C206464203100000000696C6D6300005D3E616D633C6C650000;
defparam sp_inst_23.INIT_RAM_3E = 256'h726F7373646479666F6D005D756C3C2064642034000000007479737364647966;
defparam sp_inst_23.INIT_RAM_3F = 256'h697400005D7474206D6900007465005D756F0000637500003176005D00000000;

SP sp_inst_24 (
    .DO({sp_inst_24_dout_w[15:0],sp_inst_24_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_8}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_24.READ_MODE = 1'b0;
defparam sp_inst_24.WRITE_MODE = 2'b01;
defparam sp_inst_24.BIT_WIDTH = 16;
defparam sp_inst_24.BLK_SEL = 3'b001;
defparam sp_inst_24.RESET_MODE = "SYNC";
defparam sp_inst_24.INIT_RAM_00 = 256'h20706B610000656B00005D7474206C650000616C0000747320726974726F0072;
defparam sp_inst_24.INIT_RAM_01 = 256'h6373703C63320000706300007365676400670000736563740000657400007473;
defparam sp_inst_24.INIT_RAM_02 = 256'h74613C20646465723E726170633C633200007763000061637270326900003E65;
defparam sp_inst_24.INIT_RAM_03 = 256'h000065723269005D646465723E726170633C633200007263006572773269005D;
defparam sp_inst_24.INIT_RAM_04 = 256'h3E3D616C69700000797000005D3E207474610000647400006461000063640063;
defparam sp_inst_24.INIT_RAM_05 = 256'h6E6972610000696E00003E6E746561620000706F00006172797000006873665F;
defparam sp_inst_24.INIT_RAM_06 = 256'h005D6972697000007277005D61726970006572650000696E697000006E69005D;
defparam sp_inst_24.INIT_RAM_07 = 256'h0000000074780000746E6F69005D616C69700000616C00006165697000006472;
defparam sp_inst_24.INIT_RAM_08 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C0000004C5500004C4C;
defparam sp_inst_24.INIT_RAM_09 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_24.INIT_RAM_0A = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_24.INIT_RAM_0B = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_24.INIT_RAM_0C = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_24.INIT_RAM_0D = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_24.INIT_RAM_0E = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_24.INIT_RAM_0F = 256'h00000A0A646E6D6F1C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_24.INIT_RAM_10 = 256'h3A657375000021216E616F636E69646E3A525245000A09737325000073253225;
defparam sp_inst_24.INIT_RAM_11 = 256'h6425206D00006425206E000A25203072000044430000002000003E643C206C65;
defparam sp_inst_24.INIT_RAM_12 = 256'h3A6573750000323000007838783000000D0A756E203E646120313A6573750000;
defparam sp_inst_24.INIT_RAM_13 = 256'h756C3C20646420313A6573750000383000003A78257800003E6D3C2064642034;
defparam sp_inst_24.INIT_RAM_14 = 256'h00002E2E626D2078206C656C00000D0A756C3C20646420343A65737500000D0A;
defparam sp_inst_24.INIT_RAM_15 = 256'h74732064616D4D5700000A3E6E3C72643C203A65737500002E2E626D206C656C;
defparam sp_inst_24.INIT_RAM_16 = 256'h25783D20206C435F0000726F65730000646E74732064616D4D57000064656174;
defparam sp_inst_24.INIT_RAM_17 = 256'h20202020744143202020000A25783D20546C505F000A25783D2068544F5F000A;
defparam sp_inst_24.INIT_RAM_18 = 256'h2033202020203020303020202020000A257820203825203D643200000A73746E;
defparam sp_inst_24.INIT_RAM_19 = 256'h746E000064340000767300000A31202020203020383020372020202030203430;
defparam sp_inst_24.INIT_RAM_1A = 256'h6F5400006E610000746920686F54002E745F6F64746920686F7400007469006C;
defparam sp_inst_24.INIT_RAM_1B = 256'h6E613C20745F6F646E7720686F7400006E7720686F5400006E7700006E612068;
defparam sp_inst_24.INIT_RAM_1C = 256'h203A617300006F7220746E490000776F00006C6C20686F5400006C6C00003E6C;
defparam sp_inst_24.INIT_RAM_1D = 256'h20096C656168203E5F6E643C776F6863742020200A093E686E773C206E696375;
defparam sp_inst_24.INIT_RAM_1E = 256'h7320756F2020202009206F70637520202020090961636863742020200A202020;
defparam sp_inst_24.INIT_RAM_1F = 256'h7472733C636969723C2070686567552000000A2E2E747473656D207468200077;
defparam sp_inst_24.INIT_RAM_20 = 256'h733C656D616C65675520000A3A63612E2E747473656D20656320000065733E73;
defparam sp_inst_24.INIT_RAM_21 = 256'h0000642500006425000061763E732C73322C3A31646F2079656465675520003E;
defparam sp_inst_24.INIT_RAM_22 = 256'h657370756177656755200000642567722E2E72612070656B2072695400006425;
defparam sp_inst_24.INIT_RAM_23 = 256'h00000A0D656D20797073206F65740000000021726D75666F676E206772770000;
defparam sp_inst_24.INIT_RAM_24 = 256'h3A6D6868642D2069657400000A0D6D6974656F74733A3A6864646D2D20736574;
defparam sp_inst_24.INIT_RAM_25 = 256'h74656F7465676E6969206E65726675703A202066657400000A0D6E6965737420;
defparam sp_inst_24.INIT_RAM_26 = 256'h2065646C6873000061722064617600000D72656D6170636500000A0D6C616572;
defparam sp_inst_24.INIT_RAM_27 = 256'h6432000064322D64252D3025000A6761207220686574000A482037326F74736F;
defparam sp_inst_24.INIT_RAM_28 = 256'h2E2E74727320657464771C001C001C001C000000000000000000000030253230;
defparam sp_inst_24.INIT_RAM_29 = 256'h646465723E726170633C63323A657375003E733C64776567552000000A646367;
defparam sp_inst_24.INIT_RAM_2A = 256'h61673C3E6461686363323A657375000025787264000078307461000A74613C20;
defparam sp_inst_24.INIT_RAM_2B = 256'h2820657300007365743C7669203E733C444100000D7825786174722000003E72;
defparam sp_inst_24.INIT_RAM_2C = 256'h202C7276302E352854555629202C2E312820414329322C314344312830494441;
defparam sp_inst_24.INIT_RAM_2D = 256'h3A657375000025656C75616300343A313264302069640000616329372C667629;
defparam sp_inst_24.INIT_RAM_2E = 256'h000000006574617220677277000A495032204F49203130494441203E20747461;
defparam sp_inst_24.INIT_RAM_2F = 256'h206572773A657375000A2578646900003E323C206E693A657375000A72727970;
defparam sp_inst_24.INIT_RAM_30 = 256'h6572000A72643C2065723A65737500000000000072612065727700000A206464;
defparam sp_inst_24.INIT_RAM_31 = 256'h6464206572653A657375000A3D726169253D6164726F65206568000074727320;
defparam sp_inst_24.INIT_RAM_32 = 256'h6F6B6863000A6F646172727000007261206D676F000072612065726500000A20;
defparam sp_inst_24.INIT_RAM_33 = 256'h782525207272797000007472732072696F630000656E206B6863000074727320;
defparam sp_inst_24.INIT_RAM_34 = 256'h2E2E495F4F532E2E2E2E2E2E00000A0D20203A636620203A696C3C2000000A78;
defparam sp_inst_24.INIT_RAM_35 = 256'h41422E2E2E2E2E2E000078253A6C6E617965746E63752D2D00002E2E2E2E2E2E;
defparam sp_inst_24.INIT_RAM_36 = 256'h657200000A2E2E2E2E2E2E2E44412E2E2E2E2E2E00002E2E2E2E2E2E2E2E4146;
defparam sp_inst_24.INIT_RAM_37 = 256'h1C001C001C001C001C001C001C001C001C0000002E2E7572746E726163206D69;
defparam sp_inst_24.INIT_RAM_38 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_24.INIT_RAM_39 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_24.INIT_RAM_3A = 256'h697069740072646E5F715F30697069741C001C001C001C001C001C001C001C00;
defparam sp_inst_24.INIT_RAM_3B = 256'h0072646E5F715F33697069740072646E5F715F32697069740072646E5F715F31;
defparam sp_inst_24.INIT_RAM_3C = 256'h5F715F36697069740072646E5F715F35697069740072646E5F715F3469706974;
defparam sp_inst_24.INIT_RAM_3D = 256'h697069740072646E5F715F30697069740072646E5F715F37697069740072646E;
defparam sp_inst_24.INIT_RAM_3E = 256'h0072646E5F715F33697069740072646E5F715F32697069740072646E5F715F31;
defparam sp_inst_24.INIT_RAM_3F = 256'h5F715F36697069740072646E5F715F35697069740072646E5F715F3469706974;

SP sp_inst_25 (
    .DO({sp_inst_25_dout_w[15:0],sp_inst_25_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_9}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_25.READ_MODE = 1'b0;
defparam sp_inst_25.WRITE_MODE = 2'b01;
defparam sp_inst_25.BIT_WIDTH = 16;
defparam sp_inst_25.BLK_SEL = 3'b001;
defparam sp_inst_25.RESET_MODE = "SYNC";
defparam sp_inst_25.INIT_RAM_00 = 256'h697069740072646E5F715F30697069740072646E5F715F37697069740072646E;
defparam sp_inst_25.INIT_RAM_01 = 256'h0072646E5F715F33697069740072646E5F715F32697069740072646E5F715F31;
defparam sp_inst_25.INIT_RAM_02 = 256'h5F715F36697069740072646E5F715F35697069740072646E5F715F3469706974;
defparam sp_inst_25.INIT_RAM_03 = 256'h697069740072646E5F715F30697069740072646E5F715F37697069740072646E;
defparam sp_inst_25.INIT_RAM_04 = 256'h0072646E5F715F33697069740072646E5F715F32697069740072646E5F715F31;
defparam sp_inst_25.INIT_RAM_05 = 256'h5F715F36697069740072646E5F715F35697069740072646E5F715F3469706974;
defparam sp_inst_25.INIT_RAM_06 = 256'h000000001C001C0000000072646E5F740072646E5F715F37697069740072646E;
defparam sp_inst_25.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_26 (
    .DO({sp_inst_26_dout_w[15:0],sp_inst_26_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_10}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_26.READ_MODE = 1'b0;
defparam sp_inst_26.WRITE_MODE = 2'b01;
defparam sp_inst_26.BIT_WIDTH = 16;
defparam sp_inst_26.BLK_SEL = 3'b001;
defparam sp_inst_26.RESET_MODE = "SYNC";
defparam sp_inst_26.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_27 (
    .DO({sp_inst_27_dout_w[15:0],sp_inst_27_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_11}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_27.READ_MODE = 1'b0;
defparam sp_inst_27.WRITE_MODE = 2'b01;
defparam sp_inst_27.BIT_WIDTH = 16;
defparam sp_inst_27.BLK_SEL = 3'b001;
defparam sp_inst_27.RESET_MODE = "SYNC";
defparam sp_inst_27.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_28 (
    .DO({sp_inst_28_dout_w[15:0],sp_inst_28_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_12}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_28.READ_MODE = 1'b0;
defparam sp_inst_28.WRITE_MODE = 2'b01;
defparam sp_inst_28.BIT_WIDTH = 16;
defparam sp_inst_28.BLK_SEL = 3'b001;
defparam sp_inst_28.RESET_MODE = "SYNC";
defparam sp_inst_28.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_29 (
    .DO({sp_inst_29_dout_w[15:0],sp_inst_29_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_13}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_29.READ_MODE = 1'b0;
defparam sp_inst_29.WRITE_MODE = 2'b01;
defparam sp_inst_29.BIT_WIDTH = 16;
defparam sp_inst_29.BLK_SEL = 3'b001;
defparam sp_inst_29.RESET_MODE = "SYNC";
defparam sp_inst_29.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_30 (
    .DO({sp_inst_30_dout_w[15:0],sp_inst_30_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_14}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_30.READ_MODE = 1'b0;
defparam sp_inst_30.WRITE_MODE = 2'b01;
defparam sp_inst_30.BIT_WIDTH = 16;
defparam sp_inst_30.BLK_SEL = 3'b001;
defparam sp_inst_30.RESET_MODE = "SYNC";
defparam sp_inst_30.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_31 (
    .DO({sp_inst_31_dout_w[15:0],sp_inst_31_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_15}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_31.READ_MODE = 1'b0;
defparam sp_inst_31.WRITE_MODE = 2'b01;
defparam sp_inst_31.BIT_WIDTH = 16;
defparam sp_inst_31.BLK_SEL = 3'b001;
defparam sp_inst_31.RESET_MODE = "SYNC";
defparam sp_inst_31.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
DFFRE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
DFFRE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
DFFRE dff_inst_3 (
  .Q(dff_q_3),
  .D(ad[10]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(sp_inst_0_dout[0]),
  .I1(sp_inst_1_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(sp_inst_2_dout[0]),
  .I1(sp_inst_3_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(sp_inst_4_dout[0]),
  .I1(sp_inst_5_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(sp_inst_6_dout[0]),
  .I1(sp_inst_7_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(sp_inst_8_dout[0]),
  .I1(sp_inst_9_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(sp_inst_10_dout[0]),
  .I1(sp_inst_11_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(sp_inst_12_dout[0]),
  .I1(sp_inst_13_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(sp_inst_14_dout[0]),
  .I1(sp_inst_15_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_2)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_2)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_2)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(dff_q_2)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(dff_q_1)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_1)
);
MUX2 mux_inst_14 (
  .O(dout[0]),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_0)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(sp_inst_0_dout[1]),
  .I1(sp_inst_1_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(sp_inst_2_dout[1]),
  .I1(sp_inst_3_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(sp_inst_4_dout[1]),
  .I1(sp_inst_5_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(sp_inst_6_dout[1]),
  .I1(sp_inst_7_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(sp_inst_8_dout[1]),
  .I1(sp_inst_9_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(sp_inst_10_dout[1]),
  .I1(sp_inst_11_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(sp_inst_12_dout[1]),
  .I1(sp_inst_13_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(sp_inst_14_dout[1]),
  .I1(sp_inst_15_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(mux_o_15),
  .I1(mux_o_16),
  .S0(dff_q_2)
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(mux_o_17),
  .I1(mux_o_18),
  .S0(dff_q_2)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(mux_o_19),
  .I1(mux_o_20),
  .S0(dff_q_2)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(mux_o_21),
  .I1(mux_o_22),
  .S0(dff_q_2)
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(mux_o_23),
  .I1(mux_o_24),
  .S0(dff_q_1)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(mux_o_25),
  .I1(mux_o_26),
  .S0(dff_q_1)
);
MUX2 mux_inst_29 (
  .O(dout[1]),
  .I0(mux_o_27),
  .I1(mux_o_28),
  .S0(dff_q_0)
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(sp_inst_0_dout[2]),
  .I1(sp_inst_1_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(sp_inst_2_dout[2]),
  .I1(sp_inst_3_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(sp_inst_4_dout[2]),
  .I1(sp_inst_5_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(sp_inst_6_dout[2]),
  .I1(sp_inst_7_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(sp_inst_8_dout[2]),
  .I1(sp_inst_9_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(sp_inst_10_dout[2]),
  .I1(sp_inst_11_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(sp_inst_12_dout[2]),
  .I1(sp_inst_13_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(sp_inst_14_dout[2]),
  .I1(sp_inst_15_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(dff_q_2)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(dff_q_2)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_34),
  .I1(mux_o_35),
  .S0(dff_q_2)
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(mux_o_36),
  .I1(mux_o_37),
  .S0(dff_q_2)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(dff_q_1)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(dff_q_1)
);
MUX2 mux_inst_44 (
  .O(dout[2]),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(dff_q_0)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(sp_inst_0_dout[3]),
  .I1(sp_inst_1_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(sp_inst_2_dout[3]),
  .I1(sp_inst_3_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(sp_inst_4_dout[3]),
  .I1(sp_inst_5_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(sp_inst_6_dout[3]),
  .I1(sp_inst_7_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(sp_inst_8_dout[3]),
  .I1(sp_inst_9_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(sp_inst_10_dout[3]),
  .I1(sp_inst_11_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(sp_inst_12_dout[3]),
  .I1(sp_inst_13_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(sp_inst_14_dout[3]),
  .I1(sp_inst_15_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(dff_q_2)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_47),
  .I1(mux_o_48),
  .S0(dff_q_2)
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(dff_q_2)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(mux_o_51),
  .I1(mux_o_52),
  .S0(dff_q_2)
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(mux_o_53),
  .I1(mux_o_54),
  .S0(dff_q_1)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(mux_o_55),
  .I1(mux_o_56),
  .S0(dff_q_1)
);
MUX2 mux_inst_59 (
  .O(dout[3]),
  .I0(mux_o_57),
  .I1(mux_o_58),
  .S0(dff_q_0)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(sp_inst_0_dout[4]),
  .I1(sp_inst_1_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(sp_inst_2_dout[4]),
  .I1(sp_inst_3_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(sp_inst_4_dout[4]),
  .I1(sp_inst_5_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(sp_inst_6_dout[4]),
  .I1(sp_inst_7_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(sp_inst_8_dout[4]),
  .I1(sp_inst_9_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(sp_inst_10_dout[4]),
  .I1(sp_inst_11_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(sp_inst_12_dout[4]),
  .I1(sp_inst_13_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(sp_inst_14_dout[4]),
  .I1(sp_inst_15_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(dff_q_2)
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(dff_q_2)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(mux_o_64),
  .I1(mux_o_65),
  .S0(dff_q_2)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(dff_q_2)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(mux_o_68),
  .I1(mux_o_69),
  .S0(dff_q_1)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(dff_q_1)
);
MUX2 mux_inst_74 (
  .O(dout[4]),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(dff_q_0)
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(sp_inst_0_dout[5]),
  .I1(sp_inst_1_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(sp_inst_2_dout[5]),
  .I1(sp_inst_3_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(sp_inst_4_dout[5]),
  .I1(sp_inst_5_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(sp_inst_6_dout[5]),
  .I1(sp_inst_7_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(sp_inst_8_dout[5]),
  .I1(sp_inst_9_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(sp_inst_10_dout[5]),
  .I1(sp_inst_11_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(sp_inst_12_dout[5]),
  .I1(sp_inst_13_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(sp_inst_14_dout[5]),
  .I1(sp_inst_15_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(mux_o_75),
  .I1(mux_o_76),
  .S0(dff_q_2)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(dff_q_2)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(dff_q_2)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(dff_q_2)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(mux_o_83),
  .I1(mux_o_84),
  .S0(dff_q_1)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(dff_q_1)
);
MUX2 mux_inst_89 (
  .O(dout[5]),
  .I0(mux_o_87),
  .I1(mux_o_88),
  .S0(dff_q_0)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(sp_inst_0_dout[6]),
  .I1(sp_inst_1_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(sp_inst_2_dout[6]),
  .I1(sp_inst_3_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(sp_inst_4_dout[6]),
  .I1(sp_inst_5_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(sp_inst_6_dout[6]),
  .I1(sp_inst_7_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(sp_inst_8_dout[6]),
  .I1(sp_inst_9_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(sp_inst_10_dout[6]),
  .I1(sp_inst_11_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(sp_inst_12_dout[6]),
  .I1(sp_inst_13_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(sp_inst_14_dout[6]),
  .I1(sp_inst_15_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(dff_q_2)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(dff_q_2)
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(mux_o_94),
  .I1(mux_o_95),
  .S0(dff_q_2)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_96),
  .I1(mux_o_97),
  .S0(dff_q_2)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_98),
  .I1(mux_o_99),
  .S0(dff_q_1)
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(mux_o_100),
  .I1(mux_o_101),
  .S0(dff_q_1)
);
MUX2 mux_inst_104 (
  .O(dout[6]),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(dff_q_0)
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(sp_inst_0_dout[7]),
  .I1(sp_inst_1_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(sp_inst_2_dout[7]),
  .I1(sp_inst_3_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(sp_inst_4_dout[7]),
  .I1(sp_inst_5_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(sp_inst_6_dout[7]),
  .I1(sp_inst_7_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(sp_inst_8_dout[7]),
  .I1(sp_inst_9_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(sp_inst_10_dout[7]),
  .I1(sp_inst_11_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(sp_inst_12_dout[7]),
  .I1(sp_inst_13_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(sp_inst_14_dout[7]),
  .I1(sp_inst_15_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(dff_q_2)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(dff_q_2)
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(dff_q_2)
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_111),
  .I1(mux_o_112),
  .S0(dff_q_2)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_113),
  .I1(mux_o_114),
  .S0(dff_q_1)
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_115),
  .I1(mux_o_116),
  .S0(dff_q_1)
);
MUX2 mux_inst_119 (
  .O(dout[7]),
  .I0(mux_o_117),
  .I1(mux_o_118),
  .S0(dff_q_0)
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(sp_inst_0_dout[8]),
  .I1(sp_inst_1_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(sp_inst_2_dout[8]),
  .I1(sp_inst_3_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(sp_inst_4_dout[8]),
  .I1(sp_inst_5_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(sp_inst_6_dout[8]),
  .I1(sp_inst_7_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(sp_inst_8_dout[8]),
  .I1(sp_inst_9_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_125 (
  .O(mux_o_125),
  .I0(sp_inst_10_dout[8]),
  .I1(sp_inst_11_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(sp_inst_12_dout[8]),
  .I1(sp_inst_13_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(sp_inst_14_dout[8]),
  .I1(sp_inst_15_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(mux_o_120),
  .I1(mux_o_121),
  .S0(dff_q_2)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(mux_o_122),
  .I1(mux_o_123),
  .S0(dff_q_2)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(mux_o_124),
  .I1(mux_o_125),
  .S0(dff_q_2)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(dff_q_2)
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(dff_q_1)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(dff_q_1)
);
MUX2 mux_inst_134 (
  .O(dout[8]),
  .I0(mux_o_132),
  .I1(mux_o_133),
  .S0(dff_q_0)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(sp_inst_0_dout[9]),
  .I1(sp_inst_1_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(sp_inst_2_dout[9]),
  .I1(sp_inst_3_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(sp_inst_4_dout[9]),
  .I1(sp_inst_5_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(sp_inst_6_dout[9]),
  .I1(sp_inst_7_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(sp_inst_8_dout[9]),
  .I1(sp_inst_9_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(sp_inst_10_dout[9]),
  .I1(sp_inst_11_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(sp_inst_12_dout[9]),
  .I1(sp_inst_13_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(sp_inst_14_dout[9]),
  .I1(sp_inst_15_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(mux_o_135),
  .I1(mux_o_136),
  .S0(dff_q_2)
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(dff_q_2)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(mux_o_139),
  .I1(mux_o_140),
  .S0(dff_q_2)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(mux_o_141),
  .I1(mux_o_142),
  .S0(dff_q_2)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(mux_o_143),
  .I1(mux_o_144),
  .S0(dff_q_1)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(mux_o_145),
  .I1(mux_o_146),
  .S0(dff_q_1)
);
MUX2 mux_inst_149 (
  .O(dout[9]),
  .I0(mux_o_147),
  .I1(mux_o_148),
  .S0(dff_q_0)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(sp_inst_0_dout[10]),
  .I1(sp_inst_1_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(sp_inst_2_dout[10]),
  .I1(sp_inst_3_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(sp_inst_4_dout[10]),
  .I1(sp_inst_5_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(sp_inst_6_dout[10]),
  .I1(sp_inst_7_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(sp_inst_8_dout[10]),
  .I1(sp_inst_9_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(sp_inst_10_dout[10]),
  .I1(sp_inst_11_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(sp_inst_12_dout[10]),
  .I1(sp_inst_13_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(sp_inst_14_dout[10]),
  .I1(sp_inst_15_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(mux_o_150),
  .I1(mux_o_151),
  .S0(dff_q_2)
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(mux_o_152),
  .I1(mux_o_153),
  .S0(dff_q_2)
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(mux_o_154),
  .I1(mux_o_155),
  .S0(dff_q_2)
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(mux_o_156),
  .I1(mux_o_157),
  .S0(dff_q_2)
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(mux_o_158),
  .I1(mux_o_159),
  .S0(dff_q_1)
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(mux_o_160),
  .I1(mux_o_161),
  .S0(dff_q_1)
);
MUX2 mux_inst_164 (
  .O(dout[10]),
  .I0(mux_o_162),
  .I1(mux_o_163),
  .S0(dff_q_0)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(sp_inst_0_dout[11]),
  .I1(sp_inst_1_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(sp_inst_2_dout[11]),
  .I1(sp_inst_3_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(sp_inst_4_dout[11]),
  .I1(sp_inst_5_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(sp_inst_6_dout[11]),
  .I1(sp_inst_7_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(sp_inst_8_dout[11]),
  .I1(sp_inst_9_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(sp_inst_10_dout[11]),
  .I1(sp_inst_11_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(sp_inst_12_dout[11]),
  .I1(sp_inst_13_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(sp_inst_14_dout[11]),
  .I1(sp_inst_15_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(dff_q_2)
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(mux_o_167),
  .I1(mux_o_168),
  .S0(dff_q_2)
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(mux_o_169),
  .I1(mux_o_170),
  .S0(dff_q_2)
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(mux_o_171),
  .I1(mux_o_172),
  .S0(dff_q_2)
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(mux_o_173),
  .I1(mux_o_174),
  .S0(dff_q_1)
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(mux_o_175),
  .I1(mux_o_176),
  .S0(dff_q_1)
);
MUX2 mux_inst_179 (
  .O(dout[11]),
  .I0(mux_o_177),
  .I1(mux_o_178),
  .S0(dff_q_0)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(sp_inst_0_dout[12]),
  .I1(sp_inst_1_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(sp_inst_2_dout[12]),
  .I1(sp_inst_3_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(sp_inst_4_dout[12]),
  .I1(sp_inst_5_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(sp_inst_6_dout[12]),
  .I1(sp_inst_7_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(sp_inst_8_dout[12]),
  .I1(sp_inst_9_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(sp_inst_10_dout[12]),
  .I1(sp_inst_11_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(sp_inst_12_dout[12]),
  .I1(sp_inst_13_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(sp_inst_14_dout[12]),
  .I1(sp_inst_15_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(mux_o_180),
  .I1(mux_o_181),
  .S0(dff_q_2)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(mux_o_182),
  .I1(mux_o_183),
  .S0(dff_q_2)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(mux_o_184),
  .I1(mux_o_185),
  .S0(dff_q_2)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(dff_q_2)
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(mux_o_188),
  .I1(mux_o_189),
  .S0(dff_q_1)
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(mux_o_190),
  .I1(mux_o_191),
  .S0(dff_q_1)
);
MUX2 mux_inst_194 (
  .O(dout[12]),
  .I0(mux_o_192),
  .I1(mux_o_193),
  .S0(dff_q_0)
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(sp_inst_0_dout[13]),
  .I1(sp_inst_1_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(sp_inst_2_dout[13]),
  .I1(sp_inst_3_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(sp_inst_4_dout[13]),
  .I1(sp_inst_5_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(sp_inst_6_dout[13]),
  .I1(sp_inst_7_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(sp_inst_8_dout[13]),
  .I1(sp_inst_9_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(sp_inst_10_dout[13]),
  .I1(sp_inst_11_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(sp_inst_12_dout[13]),
  .I1(sp_inst_13_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(sp_inst_14_dout[13]),
  .I1(sp_inst_15_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_195),
  .I1(mux_o_196),
  .S0(dff_q_2)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(mux_o_197),
  .I1(mux_o_198),
  .S0(dff_q_2)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_199),
  .I1(mux_o_200),
  .S0(dff_q_2)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_201),
  .I1(mux_o_202),
  .S0(dff_q_2)
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(mux_o_203),
  .I1(mux_o_204),
  .S0(dff_q_1)
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(dff_q_1)
);
MUX2 mux_inst_209 (
  .O(dout[13]),
  .I0(mux_o_207),
  .I1(mux_o_208),
  .S0(dff_q_0)
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(sp_inst_0_dout[14]),
  .I1(sp_inst_1_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(sp_inst_2_dout[14]),
  .I1(sp_inst_3_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(sp_inst_4_dout[14]),
  .I1(sp_inst_5_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(sp_inst_6_dout[14]),
  .I1(sp_inst_7_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(sp_inst_8_dout[14]),
  .I1(sp_inst_9_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(sp_inst_10_dout[14]),
  .I1(sp_inst_11_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(sp_inst_12_dout[14]),
  .I1(sp_inst_13_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(sp_inst_14_dout[14]),
  .I1(sp_inst_15_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(mux_o_210),
  .I1(mux_o_211),
  .S0(dff_q_2)
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(mux_o_212),
  .I1(mux_o_213),
  .S0(dff_q_2)
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(mux_o_214),
  .I1(mux_o_215),
  .S0(dff_q_2)
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(mux_o_216),
  .I1(mux_o_217),
  .S0(dff_q_2)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(mux_o_218),
  .I1(mux_o_219),
  .S0(dff_q_1)
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(mux_o_220),
  .I1(mux_o_221),
  .S0(dff_q_1)
);
MUX2 mux_inst_224 (
  .O(dout[14]),
  .I0(mux_o_222),
  .I1(mux_o_223),
  .S0(dff_q_0)
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(sp_inst_0_dout[15]),
  .I1(sp_inst_1_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(sp_inst_2_dout[15]),
  .I1(sp_inst_3_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(sp_inst_4_dout[15]),
  .I1(sp_inst_5_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(sp_inst_6_dout[15]),
  .I1(sp_inst_7_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(sp_inst_8_dout[15]),
  .I1(sp_inst_9_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(sp_inst_10_dout[15]),
  .I1(sp_inst_11_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(sp_inst_12_dout[15]),
  .I1(sp_inst_13_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(sp_inst_14_dout[15]),
  .I1(sp_inst_15_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_225),
  .I1(mux_o_226),
  .S0(dff_q_2)
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(mux_o_227),
  .I1(mux_o_228),
  .S0(dff_q_2)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_229),
  .I1(mux_o_230),
  .S0(dff_q_2)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(dff_q_2)
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(dff_q_1)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_1)
);
MUX2 mux_inst_239 (
  .O(dout[15]),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(dff_q_0)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(sp_inst_16_dout[16]),
  .I1(sp_inst_17_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(sp_inst_18_dout[16]),
  .I1(sp_inst_19_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(sp_inst_20_dout[16]),
  .I1(sp_inst_21_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(sp_inst_22_dout[16]),
  .I1(sp_inst_23_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(sp_inst_24_dout[16]),
  .I1(sp_inst_25_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(sp_inst_26_dout[16]),
  .I1(sp_inst_27_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(sp_inst_28_dout[16]),
  .I1(sp_inst_29_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(sp_inst_30_dout[16]),
  .I1(sp_inst_31_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(mux_o_240),
  .I1(mux_o_241),
  .S0(dff_q_2)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_242),
  .I1(mux_o_243),
  .S0(dff_q_2)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_244),
  .I1(mux_o_245),
  .S0(dff_q_2)
);
MUX2 mux_inst_251 (
  .O(mux_o_251),
  .I0(mux_o_246),
  .I1(mux_o_247),
  .S0(dff_q_2)
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(mux_o_248),
  .I1(mux_o_249),
  .S0(dff_q_1)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(mux_o_250),
  .I1(mux_o_251),
  .S0(dff_q_1)
);
MUX2 mux_inst_254 (
  .O(dout[16]),
  .I0(mux_o_252),
  .I1(mux_o_253),
  .S0(dff_q_0)
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(sp_inst_16_dout[17]),
  .I1(sp_inst_17_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(sp_inst_18_dout[17]),
  .I1(sp_inst_19_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(sp_inst_20_dout[17]),
  .I1(sp_inst_21_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(sp_inst_22_dout[17]),
  .I1(sp_inst_23_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(sp_inst_24_dout[17]),
  .I1(sp_inst_25_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(sp_inst_26_dout[17]),
  .I1(sp_inst_27_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(sp_inst_28_dout[17]),
  .I1(sp_inst_29_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(sp_inst_30_dout[17]),
  .I1(sp_inst_31_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(mux_o_255),
  .I1(mux_o_256),
  .S0(dff_q_2)
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(mux_o_257),
  .I1(mux_o_258),
  .S0(dff_q_2)
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(mux_o_259),
  .I1(mux_o_260),
  .S0(dff_q_2)
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(mux_o_261),
  .I1(mux_o_262),
  .S0(dff_q_2)
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(mux_o_263),
  .I1(mux_o_264),
  .S0(dff_q_1)
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(mux_o_265),
  .I1(mux_o_266),
  .S0(dff_q_1)
);
MUX2 mux_inst_269 (
  .O(dout[17]),
  .I0(mux_o_267),
  .I1(mux_o_268),
  .S0(dff_q_0)
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(sp_inst_16_dout[18]),
  .I1(sp_inst_17_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(sp_inst_18_dout[18]),
  .I1(sp_inst_19_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_272 (
  .O(mux_o_272),
  .I0(sp_inst_20_dout[18]),
  .I1(sp_inst_21_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(sp_inst_22_dout[18]),
  .I1(sp_inst_23_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(sp_inst_24_dout[18]),
  .I1(sp_inst_25_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(sp_inst_26_dout[18]),
  .I1(sp_inst_27_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(sp_inst_28_dout[18]),
  .I1(sp_inst_29_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(sp_inst_30_dout[18]),
  .I1(sp_inst_31_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(dff_q_2)
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(mux_o_272),
  .I1(mux_o_273),
  .S0(dff_q_2)
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(mux_o_274),
  .I1(mux_o_275),
  .S0(dff_q_2)
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(mux_o_276),
  .I1(mux_o_277),
  .S0(dff_q_2)
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(mux_o_278),
  .I1(mux_o_279),
  .S0(dff_q_1)
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(mux_o_280),
  .I1(mux_o_281),
  .S0(dff_q_1)
);
MUX2 mux_inst_284 (
  .O(dout[18]),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(dff_q_0)
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(sp_inst_16_dout[19]),
  .I1(sp_inst_17_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(sp_inst_18_dout[19]),
  .I1(sp_inst_19_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(sp_inst_20_dout[19]),
  .I1(sp_inst_21_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(sp_inst_22_dout[19]),
  .I1(sp_inst_23_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(sp_inst_24_dout[19]),
  .I1(sp_inst_25_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(sp_inst_26_dout[19]),
  .I1(sp_inst_27_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(sp_inst_28_dout[19]),
  .I1(sp_inst_29_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(sp_inst_30_dout[19]),
  .I1(sp_inst_31_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(mux_o_285),
  .I1(mux_o_286),
  .S0(dff_q_2)
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(mux_o_287),
  .I1(mux_o_288),
  .S0(dff_q_2)
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(mux_o_289),
  .I1(mux_o_290),
  .S0(dff_q_2)
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(mux_o_291),
  .I1(mux_o_292),
  .S0(dff_q_2)
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(mux_o_293),
  .I1(mux_o_294),
  .S0(dff_q_1)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(mux_o_295),
  .I1(mux_o_296),
  .S0(dff_q_1)
);
MUX2 mux_inst_299 (
  .O(dout[19]),
  .I0(mux_o_297),
  .I1(mux_o_298),
  .S0(dff_q_0)
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(sp_inst_16_dout[20]),
  .I1(sp_inst_17_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(sp_inst_18_dout[20]),
  .I1(sp_inst_19_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(sp_inst_20_dout[20]),
  .I1(sp_inst_21_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(sp_inst_22_dout[20]),
  .I1(sp_inst_23_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(sp_inst_24_dout[20]),
  .I1(sp_inst_25_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(sp_inst_26_dout[20]),
  .I1(sp_inst_27_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(sp_inst_28_dout[20]),
  .I1(sp_inst_29_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(sp_inst_30_dout[20]),
  .I1(sp_inst_31_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(mux_o_300),
  .I1(mux_o_301),
  .S0(dff_q_2)
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(mux_o_302),
  .I1(mux_o_303),
  .S0(dff_q_2)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(mux_o_304),
  .I1(mux_o_305),
  .S0(dff_q_2)
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(mux_o_306),
  .I1(mux_o_307),
  .S0(dff_q_2)
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(mux_o_308),
  .I1(mux_o_309),
  .S0(dff_q_1)
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(dff_q_1)
);
MUX2 mux_inst_314 (
  .O(dout[20]),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(dff_q_0)
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(sp_inst_16_dout[21]),
  .I1(sp_inst_17_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(sp_inst_18_dout[21]),
  .I1(sp_inst_19_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(sp_inst_20_dout[21]),
  .I1(sp_inst_21_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(sp_inst_22_dout[21]),
  .I1(sp_inst_23_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(sp_inst_24_dout[21]),
  .I1(sp_inst_25_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(sp_inst_26_dout[21]),
  .I1(sp_inst_27_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(sp_inst_28_dout[21]),
  .I1(sp_inst_29_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(sp_inst_30_dout[21]),
  .I1(sp_inst_31_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(mux_o_315),
  .I1(mux_o_316),
  .S0(dff_q_2)
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(mux_o_317),
  .I1(mux_o_318),
  .S0(dff_q_2)
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(mux_o_319),
  .I1(mux_o_320),
  .S0(dff_q_2)
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(mux_o_321),
  .I1(mux_o_322),
  .S0(dff_q_2)
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(mux_o_323),
  .I1(mux_o_324),
  .S0(dff_q_1)
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(mux_o_325),
  .I1(mux_o_326),
  .S0(dff_q_1)
);
MUX2 mux_inst_329 (
  .O(dout[21]),
  .I0(mux_o_327),
  .I1(mux_o_328),
  .S0(dff_q_0)
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(sp_inst_16_dout[22]),
  .I1(sp_inst_17_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(sp_inst_18_dout[22]),
  .I1(sp_inst_19_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(sp_inst_20_dout[22]),
  .I1(sp_inst_21_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(sp_inst_22_dout[22]),
  .I1(sp_inst_23_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(sp_inst_24_dout[22]),
  .I1(sp_inst_25_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(sp_inst_26_dout[22]),
  .I1(sp_inst_27_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(sp_inst_28_dout[22]),
  .I1(sp_inst_29_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(sp_inst_30_dout[22]),
  .I1(sp_inst_31_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(mux_o_330),
  .I1(mux_o_331),
  .S0(dff_q_2)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(mux_o_332),
  .I1(mux_o_333),
  .S0(dff_q_2)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(mux_o_334),
  .I1(mux_o_335),
  .S0(dff_q_2)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(mux_o_336),
  .I1(mux_o_337),
  .S0(dff_q_2)
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(mux_o_338),
  .I1(mux_o_339),
  .S0(dff_q_1)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(mux_o_340),
  .I1(mux_o_341),
  .S0(dff_q_1)
);
MUX2 mux_inst_344 (
  .O(dout[22]),
  .I0(mux_o_342),
  .I1(mux_o_343),
  .S0(dff_q_0)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(sp_inst_16_dout[23]),
  .I1(sp_inst_17_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(sp_inst_18_dout[23]),
  .I1(sp_inst_19_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(sp_inst_20_dout[23]),
  .I1(sp_inst_21_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(sp_inst_22_dout[23]),
  .I1(sp_inst_23_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_349 (
  .O(mux_o_349),
  .I0(sp_inst_24_dout[23]),
  .I1(sp_inst_25_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(sp_inst_26_dout[23]),
  .I1(sp_inst_27_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(sp_inst_28_dout[23]),
  .I1(sp_inst_29_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(sp_inst_30_dout[23]),
  .I1(sp_inst_31_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(mux_o_345),
  .I1(mux_o_346),
  .S0(dff_q_2)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(dff_q_2)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(mux_o_349),
  .I1(mux_o_350),
  .S0(dff_q_2)
);
MUX2 mux_inst_356 (
  .O(mux_o_356),
  .I0(mux_o_351),
  .I1(mux_o_352),
  .S0(dff_q_2)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_353),
  .I1(mux_o_354),
  .S0(dff_q_1)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_355),
  .I1(mux_o_356),
  .S0(dff_q_1)
);
MUX2 mux_inst_359 (
  .O(dout[23]),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(dff_q_0)
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(sp_inst_16_dout[24]),
  .I1(sp_inst_17_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(sp_inst_18_dout[24]),
  .I1(sp_inst_19_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(sp_inst_20_dout[24]),
  .I1(sp_inst_21_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_363 (
  .O(mux_o_363),
  .I0(sp_inst_22_dout[24]),
  .I1(sp_inst_23_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(sp_inst_24_dout[24]),
  .I1(sp_inst_25_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(sp_inst_26_dout[24]),
  .I1(sp_inst_27_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(sp_inst_28_dout[24]),
  .I1(sp_inst_29_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(sp_inst_30_dout[24]),
  .I1(sp_inst_31_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(mux_o_360),
  .I1(mux_o_361),
  .S0(dff_q_2)
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(mux_o_362),
  .I1(mux_o_363),
  .S0(dff_q_2)
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(mux_o_364),
  .I1(mux_o_365),
  .S0(dff_q_2)
);
MUX2 mux_inst_371 (
  .O(mux_o_371),
  .I0(mux_o_366),
  .I1(mux_o_367),
  .S0(dff_q_2)
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(mux_o_368),
  .I1(mux_o_369),
  .S0(dff_q_1)
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(mux_o_370),
  .I1(mux_o_371),
  .S0(dff_q_1)
);
MUX2 mux_inst_374 (
  .O(dout[24]),
  .I0(mux_o_372),
  .I1(mux_o_373),
  .S0(dff_q_0)
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(sp_inst_16_dout[25]),
  .I1(sp_inst_17_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(sp_inst_18_dout[25]),
  .I1(sp_inst_19_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_377 (
  .O(mux_o_377),
  .I0(sp_inst_20_dout[25]),
  .I1(sp_inst_21_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_378 (
  .O(mux_o_378),
  .I0(sp_inst_22_dout[25]),
  .I1(sp_inst_23_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_379 (
  .O(mux_o_379),
  .I0(sp_inst_24_dout[25]),
  .I1(sp_inst_25_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_380 (
  .O(mux_o_380),
  .I0(sp_inst_26_dout[25]),
  .I1(sp_inst_27_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_381 (
  .O(mux_o_381),
  .I0(sp_inst_28_dout[25]),
  .I1(sp_inst_29_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_382 (
  .O(mux_o_382),
  .I0(sp_inst_30_dout[25]),
  .I1(sp_inst_31_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_383 (
  .O(mux_o_383),
  .I0(mux_o_375),
  .I1(mux_o_376),
  .S0(dff_q_2)
);
MUX2 mux_inst_384 (
  .O(mux_o_384),
  .I0(mux_o_377),
  .I1(mux_o_378),
  .S0(dff_q_2)
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(mux_o_379),
  .I1(mux_o_380),
  .S0(dff_q_2)
);
MUX2 mux_inst_386 (
  .O(mux_o_386),
  .I0(mux_o_381),
  .I1(mux_o_382),
  .S0(dff_q_2)
);
MUX2 mux_inst_387 (
  .O(mux_o_387),
  .I0(mux_o_383),
  .I1(mux_o_384),
  .S0(dff_q_1)
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(mux_o_385),
  .I1(mux_o_386),
  .S0(dff_q_1)
);
MUX2 mux_inst_389 (
  .O(dout[25]),
  .I0(mux_o_387),
  .I1(mux_o_388),
  .S0(dff_q_0)
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(sp_inst_16_dout[26]),
  .I1(sp_inst_17_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(sp_inst_18_dout[26]),
  .I1(sp_inst_19_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(sp_inst_20_dout[26]),
  .I1(sp_inst_21_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(sp_inst_22_dout[26]),
  .I1(sp_inst_23_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(sp_inst_24_dout[26]),
  .I1(sp_inst_25_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(sp_inst_26_dout[26]),
  .I1(sp_inst_27_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(sp_inst_28_dout[26]),
  .I1(sp_inst_29_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(sp_inst_30_dout[26]),
  .I1(sp_inst_31_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(mux_o_390),
  .I1(mux_o_391),
  .S0(dff_q_2)
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(mux_o_392),
  .I1(mux_o_393),
  .S0(dff_q_2)
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(mux_o_394),
  .I1(mux_o_395),
  .S0(dff_q_2)
);
MUX2 mux_inst_401 (
  .O(mux_o_401),
  .I0(mux_o_396),
  .I1(mux_o_397),
  .S0(dff_q_2)
);
MUX2 mux_inst_402 (
  .O(mux_o_402),
  .I0(mux_o_398),
  .I1(mux_o_399),
  .S0(dff_q_1)
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(mux_o_400),
  .I1(mux_o_401),
  .S0(dff_q_1)
);
MUX2 mux_inst_404 (
  .O(dout[26]),
  .I0(mux_o_402),
  .I1(mux_o_403),
  .S0(dff_q_0)
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(sp_inst_16_dout[27]),
  .I1(sp_inst_17_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(sp_inst_18_dout[27]),
  .I1(sp_inst_19_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(sp_inst_20_dout[27]),
  .I1(sp_inst_21_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_408 (
  .O(mux_o_408),
  .I0(sp_inst_22_dout[27]),
  .I1(sp_inst_23_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(sp_inst_24_dout[27]),
  .I1(sp_inst_25_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(sp_inst_26_dout[27]),
  .I1(sp_inst_27_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(sp_inst_28_dout[27]),
  .I1(sp_inst_29_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_412 (
  .O(mux_o_412),
  .I0(sp_inst_30_dout[27]),
  .I1(sp_inst_31_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(mux_o_405),
  .I1(mux_o_406),
  .S0(dff_q_2)
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(mux_o_407),
  .I1(mux_o_408),
  .S0(dff_q_2)
);
MUX2 mux_inst_415 (
  .O(mux_o_415),
  .I0(mux_o_409),
  .I1(mux_o_410),
  .S0(dff_q_2)
);
MUX2 mux_inst_416 (
  .O(mux_o_416),
  .I0(mux_o_411),
  .I1(mux_o_412),
  .S0(dff_q_2)
);
MUX2 mux_inst_417 (
  .O(mux_o_417),
  .I0(mux_o_413),
  .I1(mux_o_414),
  .S0(dff_q_1)
);
MUX2 mux_inst_418 (
  .O(mux_o_418),
  .I0(mux_o_415),
  .I1(mux_o_416),
  .S0(dff_q_1)
);
MUX2 mux_inst_419 (
  .O(dout[27]),
  .I0(mux_o_417),
  .I1(mux_o_418),
  .S0(dff_q_0)
);
MUX2 mux_inst_420 (
  .O(mux_o_420),
  .I0(sp_inst_16_dout[28]),
  .I1(sp_inst_17_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_421 (
  .O(mux_o_421),
  .I0(sp_inst_18_dout[28]),
  .I1(sp_inst_19_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(sp_inst_20_dout[28]),
  .I1(sp_inst_21_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(sp_inst_22_dout[28]),
  .I1(sp_inst_23_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(sp_inst_24_dout[28]),
  .I1(sp_inst_25_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(sp_inst_26_dout[28]),
  .I1(sp_inst_27_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_426 (
  .O(mux_o_426),
  .I0(sp_inst_28_dout[28]),
  .I1(sp_inst_29_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(sp_inst_30_dout[28]),
  .I1(sp_inst_31_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(mux_o_420),
  .I1(mux_o_421),
  .S0(dff_q_2)
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(mux_o_422),
  .I1(mux_o_423),
  .S0(dff_q_2)
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(mux_o_424),
  .I1(mux_o_425),
  .S0(dff_q_2)
);
MUX2 mux_inst_431 (
  .O(mux_o_431),
  .I0(mux_o_426),
  .I1(mux_o_427),
  .S0(dff_q_2)
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(mux_o_428),
  .I1(mux_o_429),
  .S0(dff_q_1)
);
MUX2 mux_inst_433 (
  .O(mux_o_433),
  .I0(mux_o_430),
  .I1(mux_o_431),
  .S0(dff_q_1)
);
MUX2 mux_inst_434 (
  .O(dout[28]),
  .I0(mux_o_432),
  .I1(mux_o_433),
  .S0(dff_q_0)
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(sp_inst_16_dout[29]),
  .I1(sp_inst_17_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(sp_inst_18_dout[29]),
  .I1(sp_inst_19_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(sp_inst_20_dout[29]),
  .I1(sp_inst_21_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(sp_inst_22_dout[29]),
  .I1(sp_inst_23_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(sp_inst_24_dout[29]),
  .I1(sp_inst_25_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_440 (
  .O(mux_o_440),
  .I0(sp_inst_26_dout[29]),
  .I1(sp_inst_27_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(sp_inst_28_dout[29]),
  .I1(sp_inst_29_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(sp_inst_30_dout[29]),
  .I1(sp_inst_31_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(mux_o_435),
  .I1(mux_o_436),
  .S0(dff_q_2)
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(mux_o_437),
  .I1(mux_o_438),
  .S0(dff_q_2)
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(mux_o_439),
  .I1(mux_o_440),
  .S0(dff_q_2)
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(mux_o_441),
  .I1(mux_o_442),
  .S0(dff_q_2)
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(mux_o_443),
  .I1(mux_o_444),
  .S0(dff_q_1)
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(mux_o_445),
  .I1(mux_o_446),
  .S0(dff_q_1)
);
MUX2 mux_inst_449 (
  .O(dout[29]),
  .I0(mux_o_447),
  .I1(mux_o_448),
  .S0(dff_q_0)
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(sp_inst_16_dout[30]),
  .I1(sp_inst_17_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(sp_inst_18_dout[30]),
  .I1(sp_inst_19_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(sp_inst_20_dout[30]),
  .I1(sp_inst_21_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_453 (
  .O(mux_o_453),
  .I0(sp_inst_22_dout[30]),
  .I1(sp_inst_23_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(sp_inst_24_dout[30]),
  .I1(sp_inst_25_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(sp_inst_26_dout[30]),
  .I1(sp_inst_27_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(sp_inst_28_dout[30]),
  .I1(sp_inst_29_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(sp_inst_30_dout[30]),
  .I1(sp_inst_31_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(mux_o_450),
  .I1(mux_o_451),
  .S0(dff_q_2)
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(mux_o_452),
  .I1(mux_o_453),
  .S0(dff_q_2)
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(mux_o_454),
  .I1(mux_o_455),
  .S0(dff_q_2)
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(mux_o_456),
  .I1(mux_o_457),
  .S0(dff_q_2)
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(mux_o_458),
  .I1(mux_o_459),
  .S0(dff_q_1)
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(mux_o_460),
  .I1(mux_o_461),
  .S0(dff_q_1)
);
MUX2 mux_inst_464 (
  .O(dout[30]),
  .I0(mux_o_462),
  .I1(mux_o_463),
  .S0(dff_q_0)
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(sp_inst_16_dout[31]),
  .I1(sp_inst_17_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(sp_inst_18_dout[31]),
  .I1(sp_inst_19_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_467 (
  .O(mux_o_467),
  .I0(sp_inst_20_dout[31]),
  .I1(sp_inst_21_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_468 (
  .O(mux_o_468),
  .I0(sp_inst_22_dout[31]),
  .I1(sp_inst_23_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_469 (
  .O(mux_o_469),
  .I0(sp_inst_24_dout[31]),
  .I1(sp_inst_25_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_470 (
  .O(mux_o_470),
  .I0(sp_inst_26_dout[31]),
  .I1(sp_inst_27_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_471 (
  .O(mux_o_471),
  .I0(sp_inst_28_dout[31]),
  .I1(sp_inst_29_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(sp_inst_30_dout[31]),
  .I1(sp_inst_31_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_473 (
  .O(mux_o_473),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(dff_q_2)
);
MUX2 mux_inst_474 (
  .O(mux_o_474),
  .I0(mux_o_467),
  .I1(mux_o_468),
  .S0(dff_q_2)
);
MUX2 mux_inst_475 (
  .O(mux_o_475),
  .I0(mux_o_469),
  .I1(mux_o_470),
  .S0(dff_q_2)
);
MUX2 mux_inst_476 (
  .O(mux_o_476),
  .I0(mux_o_471),
  .I1(mux_o_472),
  .S0(dff_q_2)
);
MUX2 mux_inst_477 (
  .O(mux_o_477),
  .I0(mux_o_473),
  .I1(mux_o_474),
  .S0(dff_q_1)
);
MUX2 mux_inst_478 (
  .O(mux_o_478),
  .I0(mux_o_475),
  .I1(mux_o_476),
  .S0(dff_q_1)
);
MUX2 mux_inst_479 (
  .O(dout[31]),
  .I0(mux_o_477),
  .I1(mux_o_478),
  .S0(dff_q_0)
);
endmodule //blk_mem_gen_0
