parameter DIN_WIDTH = 8;
parameter COEFF_WIDTH = 16;
parameter DOUT_WIDTH = 16;
parameter NUM_CHN = 1;
parameter NUM_FACTOR = 1;
parameter TAPS_SIZE = 8;
parameter NUM_TDM = 1;
parameter COEFF_PATH = "./coeff.dat";
