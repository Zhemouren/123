//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9 (64-bit)
//Part Number: GW5A-LV25MG121NES
//Device: GW5A-25
//Device Version: A
//Created Time: Fri May 17 16:22:06 2024

module Gowin_SP (dout, clk, oce, ce, reset, wre, ad, din, byte_en);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [13:0] ad;
input [31:0] din;
input [3:0] byte_en;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire [15:0] sp_inst_0_dout_w;
wire [15:0] sp_inst_0_dout;
wire [15:0] sp_inst_1_dout_w;
wire [15:0] sp_inst_1_dout;
wire [15:0] sp_inst_2_dout_w;
wire [15:0] sp_inst_2_dout;
wire [15:0] sp_inst_3_dout_w;
wire [15:0] sp_inst_3_dout;
wire [15:0] sp_inst_4_dout_w;
wire [15:0] sp_inst_4_dout;
wire [15:0] sp_inst_5_dout_w;
wire [15:0] sp_inst_5_dout;
wire [15:0] sp_inst_6_dout_w;
wire [15:0] sp_inst_6_dout;
wire [15:0] sp_inst_7_dout_w;
wire [15:0] sp_inst_7_dout;
wire [15:0] sp_inst_8_dout_w;
wire [15:0] sp_inst_8_dout;
wire [15:0] sp_inst_9_dout_w;
wire [15:0] sp_inst_9_dout;
wire [15:0] sp_inst_10_dout_w;
wire [15:0] sp_inst_10_dout;
wire [15:0] sp_inst_11_dout_w;
wire [15:0] sp_inst_11_dout;
wire [15:0] sp_inst_12_dout_w;
wire [15:0] sp_inst_12_dout;
wire [15:0] sp_inst_13_dout_w;
wire [15:0] sp_inst_13_dout;
wire [15:0] sp_inst_14_dout_w;
wire [15:0] sp_inst_14_dout;
wire [15:0] sp_inst_15_dout_w;
wire [15:0] sp_inst_15_dout;
wire [15:0] sp_inst_16_dout_w;
wire [31:16] sp_inst_16_dout;
wire [15:0] sp_inst_17_dout_w;
wire [31:16] sp_inst_17_dout;
wire [15:0] sp_inst_18_dout_w;
wire [31:16] sp_inst_18_dout;
wire [15:0] sp_inst_19_dout_w;
wire [31:16] sp_inst_19_dout;
wire [15:0] sp_inst_20_dout_w;
wire [31:16] sp_inst_20_dout;
wire [15:0] sp_inst_21_dout_w;
wire [31:16] sp_inst_21_dout;
wire [15:0] sp_inst_22_dout_w;
wire [31:16] sp_inst_22_dout;
wire [15:0] sp_inst_23_dout_w;
wire [31:16] sp_inst_23_dout;
wire [15:0] sp_inst_24_dout_w;
wire [31:16] sp_inst_24_dout;
wire [15:0] sp_inst_25_dout_w;
wire [31:16] sp_inst_25_dout;
wire [15:0] sp_inst_26_dout_w;
wire [31:16] sp_inst_26_dout;
wire [15:0] sp_inst_27_dout_w;
wire [31:16] sp_inst_27_dout;
wire [15:0] sp_inst_28_dout_w;
wire [31:16] sp_inst_28_dout;
wire [15:0] sp_inst_29_dout_w;
wire [31:16] sp_inst_29_dout;
wire [15:0] sp_inst_30_dout_w;
wire [31:16] sp_inst_30_dout;
wire [15:0] sp_inst_31_dout_w;
wire [31:16] sp_inst_31_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_60;
wire mux_o_61;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_123;
wire mux_o_124;
wire mux_o_125;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_154;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_245;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_251;
wire mux_o_252;
wire mux_o_253;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_258;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_265;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_270;
wire mux_o_271;
wire mux_o_272;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_278;
wire mux_o_279;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_308;
wire mux_o_309;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_321;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_335;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_349;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_356;
wire mux_o_357;
wire mux_o_358;
wire mux_o_360;
wire mux_o_361;
wire mux_o_362;
wire mux_o_363;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_370;
wire mux_o_371;
wire mux_o_372;
wire mux_o_373;
wire mux_o_375;
wire mux_o_376;
wire mux_o_377;
wire mux_o_378;
wire mux_o_379;
wire mux_o_380;
wire mux_o_381;
wire mux_o_382;
wire mux_o_383;
wire mux_o_384;
wire mux_o_385;
wire mux_o_386;
wire mux_o_387;
wire mux_o_388;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_401;
wire mux_o_402;
wire mux_o_403;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_408;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_412;
wire mux_o_413;
wire mux_o_414;
wire mux_o_415;
wire mux_o_416;
wire mux_o_417;
wire mux_o_418;
wire mux_o_420;
wire mux_o_421;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_426;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_431;
wire mux_o_432;
wire mux_o_433;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_440;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_453;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_460;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_465;
wire mux_o_466;
wire mux_o_467;
wire mux_o_468;
wire mux_o_469;
wire mux_o_470;
wire mux_o_471;
wire mux_o_472;
wire mux_o_473;
wire mux_o_474;
wire mux_o_475;
wire mux_o_476;
wire mux_o_477;
wire mux_o_478;
wire ce_w;
wire gw_gnd;

assign ce_w = ~wre & ce;
assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_0.INIT = 16'h0001;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_1.INIT = 16'h0002;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_2.INIT = 16'h0004;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_3.INIT = 16'h0008;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_4.INIT = 16'h0010;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_5.INIT = 16'h0020;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_6.INIT = 16'h0040;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_7.INIT = 16'h0080;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_8.INIT = 16'h0100;
LUT4 lut_inst_9 (
  .F(lut_f_9),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_9.INIT = 16'h0200;
LUT4 lut_inst_10 (
  .F(lut_f_10),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_10.INIT = 16'h0400;
LUT4 lut_inst_11 (
  .F(lut_f_11),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_11.INIT = 16'h0800;
LUT4 lut_inst_12 (
  .F(lut_f_12),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_12.INIT = 16'h1000;
LUT4 lut_inst_13 (
  .F(lut_f_13),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_13.INIT = 16'h2000;
LUT4 lut_inst_14 (
  .F(lut_f_14),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_14.INIT = 16'h4000;
LUT4 lut_inst_15 (
  .F(lut_f_15),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_15.INIT = 16'h8000;
SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[15:0],sp_inst_0_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 16;
defparam sp_inst_0.BLK_SEL = 3'b001;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h000CD1CF358E71EF002F018C002C11AD020F3590020F35F021EF018F2000000D;
defparam sp_inst_0.INIT_RAM_01 = 256'hFD8CE3EC118CFD8C002C102C000C302C002CF9AC118C018011AC51AD000D018C;
defparam sp_inst_0.INIT_RAM_02 = 256'h00000000000000000020800000203400F06300230180200C402C418CA06C442C;
defparam sp_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[15:0],sp_inst_1_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_1}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b00;
defparam sp_inst_1.BIT_WIDTH = 16;
defparam sp_inst_1.BLK_SEL = 3'b001;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'h92A8A2A7B2A6C2A5D2A472B482B392B2A2B1B2B0C2AFD2AEE2ADF2AC0055C435;
defparam sp_inst_1.INIT_RAM_01 = 256'h2DA0818D2DA0418D2DA0218D2DA0118D65A0F18D140C42A352A162AB72AA82A9;
defparam sp_inst_1.INIT_RAM_02 = 256'h140060001C00D4002400BC002C008800340004003C00C4002DA0018D2DA0018D;
defparam sp_inst_1.INIT_RAM_03 = 256'hC2A5D2A472B482B392B2A2B1B2B0C2AFD2AEE2ADF2AC0055040074000DA0018D;
defparam sp_inst_1.INIT_RAM_04 = 256'h30760000042040763076C0633800C41542A352A162AB72AA82A992A8A2A7B2A6;
defparam sp_inst_1.INIT_RAM_05 = 256'hA2C5B2C48076707680630020406330760000102C040C40763076C06300204063;
defparam sp_inst_1.INIT_RAM_06 = 256'hBECC008C80766076706180630020806370760000318DB2CC31ADA2CC318DB2CC;
defparam sp_inst_1.INIT_RAM_07 = 256'h52C662C572C4C076A076B061406300208063607670610000EC00D0040185BECC;
defparam sp_inst_1.INIT_RAM_08 = 256'h52CC5000B2C092CC72CC0C0087FFB40492CC300C72CC1D8072CC258042CC42C7;
defparam sp_inst_1.INIT_RAM_09 = 256'hB2CC92CC000709A035CC92CE52CDC1AC35CDC2CEB2CD5DCC00070980B1AE92CD;
defparam sp_inst_1.INIT_RAM_0A = 256'h1D8DB2CCA2CD7400A2CC31CC358CB5CE31ADB2CEB2CD62CCB19F92CCB2CC058C;
defparam sp_inst_1.INIT_RAM_0B = 256'h1400818CC18C818C82CC198D240C82CD82CC000C0800C18C31ACC2CDFD8CA2CC;
defparam sp_inst_1.INIT_RAM_0C = 256'hC063A076B0610184000C8C0CA2CCA2CCFD8CA2CC97FF0184818C5D8C818C82CC;
defparam sp_inst_1.INIT_RAM_0D = 256'h72CC33FF0184BECC3FFF34040DAC280CBECD300072C4C076A076B06140630020;
defparam sp_inst_1.INIT_RAM_0E = 256'hE076F06180630020C063A076B0610184000CC59FBECCBECC018C72CC72CC058C;
defparam sp_inst_1.INIT_RAM_0F = 256'h3000B2C0A2CC72CC72CC918C82CC72CB62CA52C942C832C722C612C532C40076;
defparam sp_inst_1.INIT_RAM_10 = 256'h6D8C018C31AC32CD058CB2CC92CC040CE5AC940C8ECD8ECC018C31AC32CDB2CC;
defparam sp_inst_1.INIT_RAM_11 = 256'hB2CCA2CC118CA2CCDBFF0184018CA2CC0180018C31AC118C014C898DADAC4C0D;
defparam sp_inst_1.INIT_RAM_12 = 256'hA2CC6800B2CC058CB2CCA2CC118CA2CC0FFF0184818C018CA2CC9800B2CC058C;
defparam sp_inst_1.INIT_RAM_13 = 256'h0407018CA2CC3000B2CC058CB2CCA2CC118CA2CC13FF018492C528060007018C;
defparam sp_inst_1.INIT_RAM_14 = 256'h92C520060007018CA2CCF800B2CC058CB2CCA2CC118CA2CCDBFF018492C52806;
defparam sp_inst_1.INIT_RAM_15 = 256'h6BFF018492C508060007018CA2CCC000B2CC058CB2CCA2CC118CA2CCA3FF0184;
defparam sp_inst_1.INIT_RAM_16 = 256'h118CA2CC33FF018492C540060007018CA2CC8800B2CC058CB2CCA2CC118CA2CC;
defparam sp_inst_1.INIT_RAM_17 = 256'h3C0092C0B2CC058CB2CC3800B2CC058CB2CCD3FF94045000B2CC058CB2CCA2CC;
defparam sp_inst_1.INIT_RAM_18 = 256'h058CB2CCB2CC058CB2CC92CC31AC418C018C31CC32CE058CB2CC31AD280C92CD;
defparam sp_inst_1.INIT_RAM_19 = 256'h92CD3C0092C0BBFF958DE40C018D31AC32CD058CB2CCD98DC00C018D31AC32CD;
defparam sp_inst_1.INIT_RAM_1A = 256'h32CD058CB2CCB2CC058CB2CC92CC31AC418C018C31CC32CE058CB2CC31AD280C;
defparam sp_inst_1.INIT_RAM_1B = 256'h24000000B7FF94043FFF958DE40C018D31AC32CD058CB2CC5D8DC00C018D31AC;
defparam sp_inst_1.INIT_RAM_1C = 256'hC59F018C31AC32CDB2CCB2CC058CB2CC8FFF01848ECC9BFF34040DAC280C8ECD;
defparam sp_inst_1.INIT_RAM_1D = 256'hB2CC1C00B2CC72CC52C662C572C4C076B076406300208063E076F0610184000C;
defparam sp_inst_1.INIT_RAM_1E = 256'h707680630020C063B076018472CCDD9F52CDFD8D52CC018D81AD62CDB2CD058D;
defparam sp_inst_1.INIT_RAM_1F = 256'h806370760000018DAECDB2CCF19F818C818C158CB2CC0000AECC00ACB2C48076;
defparam sp_inst_1.INIT_RAM_20 = 256'h72C4C076B07640630020406330760000D18DA9ADB4ADD60C40763076C0630020;
defparam sp_inst_1.INIT_RAM_21 = 256'hD60C018E300C31CCB2CC040E018DD60C318062CCB2CC72CC698D7C0C72CD62C5;
defparam sp_inst_1.INIT_RAM_22 = 256'hB2CC818C72CC6800018D39ADD60C018E31CCB2CC040E018DD60C9000018DB9AD;
defparam sp_inst_1.INIT_RAM_23 = 256'h040E418DD60C2800418DB9ADD60C018E300C31CCB2CC040E418DD60C318062CC;
defparam sp_inst_1.INIT_RAM_24 = 256'h72CD62C572C4C076B07640630020C063B0760000418D39ADD60C018E31CCB2CC;
defparam sp_inst_1.INIT_RAM_25 = 256'h118DB9ADD60C018E300C31CCB2CC040E118DD60C318062CCB2CC72CC698D7C0C;
defparam sp_inst_1.INIT_RAM_26 = 256'h318062CCB2CC818C72CC6800118D39ADD60C018E31CCB2CC040E118DD60C9000;
defparam sp_inst_1.INIT_RAM_27 = 256'h31CCB2CC040E518DD60C2800518DB9ADD60C018E300C31CCB2CC040E518DD60C;
defparam sp_inst_1.INIT_RAM_28 = 256'h72CC458D7C0C72CD72C4C076B07640630020C063B0760000518D39ADD60C018E;
defparam sp_inst_1.INIT_RAM_29 = 256'h72CC4400000C4C00040C0D8D35CDB2CD040EB58C35CDB2CD040E218CD60CB2CC;
defparam sp_inst_1.INIT_RAM_2A = 256'h0184000C0800040C0D8D35CDB2CD040EB58C35CDB2CD040E618CD60CB2CC818C;
defparam sp_inst_1.INIT_RAM_2B = 256'h0020806370760000F59FB2CDFD8DB2CC0000B2C48076707680630020C063B076;
defparam sp_inst_1.INIT_RAM_2C = 256'h70760000198D080DB2CC118D800DB2CC018D81AD030DB2CCB2C4807670768063;
defparam sp_inst_1.INIT_RAM_2D = 256'hB2CCB2CCA00C098D800DD20CA2CC018CD08CB2C072C4C076B076406300208063;
defparam sp_inst_1.INIT_RAM_2E = 256'h72CC098D880DD20C058D81ADD20CA18DB2CC018D81ADB2CDD20CB2CCFD8C898C;
defparam sp_inst_1.INIT_RAM_2F = 256'hD20C1580B2CCB2C48076707680630020C063B0760000118D100DD20C1180198C;
defparam sp_inst_1.INIT_RAM_30 = 256'h1580B2CCB2C48076707680630020806370760000118DFC0DD20C1000118D000D;
defparam sp_inst_1.INIT_RAM_31 = 256'h008C80766076706180630020806370760000118DFC0DD20C1000118D000DD20C;
defparam sp_inst_1.INIT_RAM_32 = 256'h80767076806300208063607670610000118D400DD20C0D8DBECDD20C7800BECC;
defparam sp_inst_1.INIT_RAM_33 = 256'h80630020806370760000ED9F098CBECCBECC118CD20C1000A2C0BECC118CD20C;
defparam sp_inst_1.INIT_RAM_34 = 256'hC0630020806370760000118D100DD20C1180118CBECCBECC118CD20C80767076;
defparam sp_inst_1.INIT_RAM_35 = 256'hD80C118D01AD006DC18CD80C018D01AD138DC18CD80C2180C18CD80C40763076;
defparam sp_inst_1.INIT_RAM_36 = 256'h31CD240C31AE000CB2CDB2C48076707680630020406330760000218D040DC18C;
defparam sp_inst_1.INIT_RAM_37 = 256'h008C8076707680630020806370760000118DC18CD80C31AD018C006C00070980;
defparam sp_inst_1.INIT_RAM_38 = 256'h8063707600000D8D81AD0DADCE0C818D898CBECC018D81AD0DADBECDCE0CBECC;
defparam sp_inst_1.INIT_RAM_39 = 256'h81AD41ADCE0C818D018CCE0C8FFF0184BECCBECC008C80766076706180630020;
defparam sp_inst_1.INIT_RAM_3A = 256'h607670610000F19F058C818C058CCE0C0000F19F118C818C058CCE0C0000018D;
defparam sp_inst_1.INIT_RAM_3B = 256'hCE0C818E158CCE0C158D81AD09ADCE0C818D158CCE0C40763076C06300208063;
defparam sp_inst_1.INIT_RAM_3C = 256'h09ADCE0C818D158CCE0C40763076C0630020406330760000158D81ADB5CD7C0D;
defparam sp_inst_1.INIT_RAM_3D = 256'h6076706180630020406330760000158D81AD81ADCE0C818D158CCE0C158D81AD;
defparam sp_inst_1.INIT_RAM_3E = 256'h80636076706100004C00C084FFC40185BECC018D040D218CFFECBECC008C8076;
defparam sp_inst_1.INIT_RAM_3F = 256'h62CCA2CCB2CC8C0072CC8580018C62CCB2CC72CC62C572C4C076B07640630020;

SP sp_inst_2 (
    .DO({sp_inst_2_dout_w[15:0],sp_inst_2_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_2}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_2.READ_MODE = 1'b0;
defparam sp_inst_2.WRITE_MODE = 2'b00;
defparam sp_inst_2.BIT_WIDTH = 16;
defparam sp_inst_2.BLK_SEL = 3'b001;
defparam sp_inst_2.RESET_MODE = "SYNC";
defparam sp_inst_2.INIT_RAM_00 = 256'h018DA2CC1980018C92CC2580018CA2CC92CC058C92CCA2CC058CA2CC1C0092CC;
defparam sp_inst_2.INIT_RAM_01 = 256'h0184000C819F018CB2CCB2CC058CB2CC2000B2CC0D80018C92CCC1AC018C92CC;
defparam sp_inst_2.INIT_RAM_02 = 256'hBECDD00CF19F818C818C158CD00C0000BECC008C8076707680630020C063B076;
defparam sp_inst_2.INIT_RAM_03 = 256'h93FFBC0467FF8084FFE400054006407620763061C0630020806370760000018D;
defparam sp_inst_2.INIT_RAM_04 = 256'h818CE18C018CC18CFFEC407620763061C063002040632076306100008BFF0404;
defparam sp_inst_2.INIT_RAM_05 = 256'h13FF0184818CA18C018CE18CFFEC2FFF0184818CC18C018C518CFFEC4BFF0184;
defparam sp_inst_2.INIT_RAM_06 = 256'h008C807660767061806300204063207630610000FBFF0184818C018C718CFFEC;
defparam sp_inst_2.INIT_RAM_07 = 256'hA18CB2CCB2C4807660767061806300208063607670610000C3FF0184BECCBECC;
defparam sp_inst_2.INIT_RAM_08 = 256'h80766076706180630020806360767061000077FF0184818CB2CC87FF0184818C;
defparam sp_inst_2.INIT_RAM_09 = 256'hBACC008C8076607670618063002080636076706100003FFF0184BECCBECC008C;
defparam sp_inst_2.INIT_RAM_0A = 256'h806300208063607670610000EBFF0184818CBACCFBFF0184818C818CA18CBACC;
defparam sp_inst_2.INIT_RAM_0B = 256'hA1ADFFED2C00A2C033FFEFFF258D040DD18CFFECB2CC418C004C807660767061;
defparam sp_inst_2.INIT_RAM_0C = 256'h058C818C158CD00C0000D18D240CA2CDA2CC058CA2CC7FFF0184018C31ACA2CC;
defparam sp_inst_2.INIT_RAM_0D = 256'h098D81AD35CDF40DD00C818E098CD00C2980B2CCB2CCFD8CB2CCA80092C0F19F;
defparam sp_inst_2.INIT_RAM_0E = 256'h018CD00C2400018031AC92CCB1ADFFED1D80B2CCB99F058C818C158CD00C1800;
defparam sp_inst_2.INIT_RAM_0F = 256'hFFEC8D8D2C0C92CD92CC058C92CCB2CCC18C00EC018D31CC92CC21CEFFEE818D;
defparam sp_inst_2.INIT_RAM_10 = 256'h0804407620763061C06300208063607670610184040C0800000C0D80258C418C;
defparam sp_inst_2.INIT_RAM_11 = 256'hB2CC3ACC3ACC008C0076E076F061006300204063207630610184008C7BFFF000;
defparam sp_inst_2.INIT_RAM_12 = 256'h7ECC818CC18C018CD18CFFEC7ACC818CE18C018C318CFFEC76CC040C72CCBC0C;
defparam sp_inst_2.INIT_RAM_13 = 256'hD00C00008EC08ACC1C0C86CC818C018C118CFFEC82CC818CA18C018C718CFFEC;
defparam sp_inst_2.INIT_RAM_14 = 256'hF40DD00C818E098CD00C2980B2CCB2CCFD8CB2CCC000A2C0F19F058C818C158C;
defparam sp_inst_2.INIT_RAM_15 = 256'h018031ACA2CC81ADFFED1D80B2CCB99F058C818C158CD00C1800098D81AD35CD;
defparam sp_inst_2.INIT_RAM_16 = 256'h2C000184018C31ACA2CCA1ADFFED018D31CCA2CCF1CEFFEE818D018CD00C2400;
defparam sp_inst_2.INIT_RAM_17 = 256'h0D8092CC92C4D7FF9084FFE4018572CC758D600CA2CDA2CC058CA2CCB2CC3ACC;
defparam sp_inst_2.INIT_RAM_18 = 256'h73FF0404EBFFA7FF807660767061806300200063E076F0610184000C080092CC;
defparam sp_inst_2.INIT_RAM_19 = 256'hA2CC1580A2CCA2C4F7FF4184004C0BFF0184B2CCB2CC140CE7FF0404A3FF0C04;
defparam sp_inst_2.INIT_RAM_1A = 256'h008CC076A076B061406300208063607670610184BECCBECCFC0C0C00BECC258C;
defparam sp_inst_2.INIT_RAM_1B = 256'hB2CC1D8C818C7ECCA3FF01847ECC53FF08040FFF1004DFFF040457FF13FF7ECC;
defparam sp_inst_2.INIT_RAM_1C = 256'hBECCBECCFC0C0C00BECC258CA2CC1580A2CCA2C44FFF4184004C63FF0184B2CC;
defparam sp_inst_2.INIT_RAM_1D = 256'h0C046FFF0C043FFF0404B7FF73FF80766076706180630020C063A076B0610184;
defparam sp_inst_2.INIT_RAM_1E = 256'h0C00BECC258CA2CC1580A2CCA2C4C3FF4184004CD7FF0184B2CCB2CC1C0CB3FF;
defparam sp_inst_2.INIT_RAM_1F = 256'hB3FF04042BFFE7FF807660767061806300208063607670610184BECCBECCFC0C;
defparam sp_inst_2.INIT_RAM_20 = 256'hA2CC1580A2CCA2C437FF4184004C4BFF0184B2CCB2CC240C27FF1404E3FF0C04;
defparam sp_inst_2.INIT_RAM_21 = 256'h008CC076A076B061406300208063607670610184BECCBECCFC0C0C00BECC258C;
defparam sp_inst_2.INIT_RAM_22 = 256'h72CCD7FF01847ECC87FF180443FF180413FF04048BFF47FF72CC01AC7ECC00AD;
defparam sp_inst_2.INIT_RAM_23 = 256'h818C818C818CA18C72CC818D7ECCAFFF0184818C72CCBFFF0184818C818CA18C;
defparam sp_inst_2.INIT_RAM_24 = 256'hA2C42BFF4184004C3FFF0184B2CCB2CC358C818C31AC818C818C72CC818D31AC;
defparam sp_inst_2.INIT_RAM_25 = 256'h706180630020C063A076B0610184BECCBECCFC0C0C00BECC258CA2CC1580A2CC;
defparam sp_inst_2.INIT_RAM_26 = 256'h004CB3FF0184B2CCB2CC440C8FFF34044BFF0C041BFF040493FF4FFF80766076;
defparam sp_inst_2.INIT_RAM_27 = 256'h8063607670610184BECCBECCFC0C0C00BECC258CA2CC1580A2CCA2C49FFF4184;
defparam sp_inst_2.INIT_RAM_28 = 256'hE3FF9FFF6ACC01AC72CC01CC7ECC52C700CD00AE008CC076A076B06140630020;
defparam sp_inst_2.INIT_RAM_29 = 256'h72CC17FF0184818C818CA18C72CC2FFF01847ECCDFFF6C049BFF20046BFF0404;
defparam sp_inst_2.INIT_RAM_2A = 256'h72CC818D7ECCDFFF0184818C6ACCEFFF0184818C818CA18C6ACC07FF0184818C;
defparam sp_inst_2.INIT_RAM_2B = 256'h818C6ACC818D31AC818CA18C6ACC818D31AC818C818C72CC818D31AC818CA18C;
defparam sp_inst_2.INIT_RAM_2C = 256'h258CA2CC8580A2CCA2C43BFF4184004C4FFF0184B2CCB2CC918C818C31AC818C;
defparam sp_inst_2.INIT_RAM_2D = 256'hA2CC018D52CC818D31AC818C018C2D8CA2CC818DA18C818C018C298CA2CCBECC;
defparam sp_inst_2.INIT_RAM_2E = 256'hBECCFC0C0C00098D52CC818D31AC818C018C358CA2CC818DA18C818C018C318C;
defparam sp_inst_2.INIT_RAM_2F = 256'h0805F80608079C007ECC008CC076A076B06140630020C063A076B0610184BECC;
defparam sp_inst_2.INIT_RAM_30 = 256'h000000000000000000008400B2CCAD8C556CC400F804080518060807D8007804;
defparam sp_inst_2.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_32 = 256'hD000759FB2CDFD8DB2CC00000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_33 = 256'h0020C063A076B0610000F40078040805E8061007B8000C006404080520061407;
defparam sp_inst_2.INIT_RAM_34 = 256'hBACC0180018C31AC218C010C898D15AC100DB6CCB2C0B6C0C076A076B0614063;
defparam sp_inst_2.INIT_RAM_35 = 256'h008C37FF040469807ECC7ECC008CC3FF800078040805E80610074400BACC058C;
defparam sp_inst_2.INIT_RAM_36 = 256'h040CBAC0280020040805340604073C00A0040805F8060807000041807ECC7ECC;
defparam sp_inst_2.INIT_RAM_37 = 256'hF80608079800BACC058CBACC5000FBFF01847ECC60000BFF01847ECC7000B6CC;
defparam sp_inst_2.INIT_RAM_38 = 256'h008C77FF080469807ECC7ECC008C03FFC0002004080534060407D400A0040805;
defparam sp_inst_2.INIT_RAM_39 = 256'h080CBAC0680020040805340604077C00A0040805F8060807400041807ECC7ECC;
defparam sp_inst_2.INIT_RAM_3A = 256'h2000A0040805F8060807E40090003BFF01847ECCA0004BFF01847ECCB000B6CC;
defparam sp_inst_2.INIT_RAM_3B = 256'hE000A0040805F8060807A40069807ECC7ECC008C83FF0C002004080534060407;
defparam sp_inst_2.INIT_RAM_3C = 256'hA000F804080508060807B40078040805F80608077800CC002004080534060407;
defparam sp_inst_2.INIT_RAM_3D = 256'h01847ECC6800F8040805100608077C0078040805F80608074000EC00B6CC0C0C;
defparam sp_inst_2.INIT_RAM_3E = 256'h000000000000000000000000000000008400A2CCC98C0E2CA800B6C0BAC05BFF;
defparam sp_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_3 (
    .DO({sp_inst_3_dout_w[15:0],sp_inst_3_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_3}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_3.READ_MODE = 1'b0;
defparam sp_inst_3.WRITE_MODE = 2'b00;
defparam sp_inst_3.BIT_WIDTH = 16;
defparam sp_inst_3.BLK_SEL = 3'b001;
defparam sp_inst_3.RESET_MODE = "SYNC";
defparam sp_inst_3.INIT_RAM_00 = 256'h7ECC7ECC008CB3FF759FA2CDFD8DA2CC00000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_01 = 256'hBECDBECC008C98009000B2CC040CD4007FFF01847ECCB6C0E800B6CC100C1180;
defparam sp_inst_3.INIT_RAM_02 = 256'hB2CC118D1C0CB2CDBEC021AC380CBECDB2CCFD8CB2CC1180B2CCBEC01DAC340C;
defparam sp_inst_3.INIT_RAM_03 = 256'hBECD2C00F0041005018604074008B2CCDC008004100580C601060807B2CC058C;
defparam sp_inst_3.INIT_RAM_04 = 256'h0805F80618075C00F5807ECC7ECC008C53FF08040185818CB2CCBEC06DAC3C0C;
defparam sp_inst_3.INIT_RAM_05 = 256'h2AACAC00F0041005018604074008B2CC5C008004100580C60106080798002804;
defparam sp_inst_3.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000840092CC598C;
defparam sp_inst_3.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_08 = 256'h82CCC98C0E2C0000AFFF01847ECCB6C0CC00759F92CDFD8D92CC000000000000;
defparam sp_inst_3.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000008400;
defparam sp_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0B = 256'hB06140630020C063A076B06100003BFF09AC280CBACD759F82CDFD8D82CC0000;
defparam sp_inst_3.INIT_RAM_0C = 256'h008C77FF0404F19F8ECC8ECC008C03FFC00078040805E80610078400C076A076;
defparam sp_inst_3.INIT_RAM_0D = 256'h7000200418006D808ECC8ECC008CA7FF040400058C06018772CC45808ECC8ECC;
defparam sp_inst_3.INIT_RAM_0E = 256'h00000000000000000000000000000000000000008400B2CCE58C472CE0008400;
defparam sp_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_10 = 256'hE58C472CB800240404003C00759FB2CDFD8DB2CC000000000000000000000000;
defparam sp_inst_3.INIT_RAM_11 = 256'h000000000000000000000000000000000000000000000000000000008400A2CC;
defparam sp_inst_3.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_13 = 256'h0000840092CC918C1C6C480008001804B000D000759FA2CDFD8DA2CC00000000;
defparam sp_inst_3.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_15 = 256'h92CC000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_16 = 256'h80630020C063A076B06100007FFF3C0078040805E80610070000759F92CDFD8D;
defparam sp_inst_3.INIT_RAM_17 = 256'hB2CC918C1C6CEBFF0184AECC100050000D80AECCAECC008CAFFF807660767061;
defparam sp_inst_3.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000008400;
defparam sp_inst_3.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1A = 256'hB2C4B2C4807660767061806300208063607670610000759FB2CDFD8DB2CC0000;
defparam sp_inst_3.INIT_RAM_1B = 256'h4063207630610000BFFF0004407620763061C06300208063607670610000DFFF;
defparam sp_inst_3.INIT_RAM_1C = 256'h407620763061C0630020406320763061000093FFBC04407620763061C0630020;
defparam sp_inst_3.INIT_RAM_1D = 256'h35CC72CD018E018CFFCC72C4C076B07640630020406320763061000067FF0004;
defparam sp_inst_3.INIT_RAM_1E = 256'h018D81ADB2CDD00C058D81ADD00CA18DB2CC0D8D000DD00CB2CCFD8C000709A0;
defparam sp_inst_3.INIT_RAM_1F = 256'h0000BECC008C8076707680630020C063B07600000D8D0C0DD00C098D180DD00C;
defparam sp_inst_3.INIT_RAM_20 = 256'h008C8076707680630020806370760000018DBECDD00CF19F818C818C158CD00C;
defparam sp_inst_3.INIT_RAM_21 = 256'h818C098CD00C098D81ADFDADD00C818D098CD00CBECC0C0C0D8D0C0CBECDBECC;
defparam sp_inst_3.INIT_RAM_22 = 256'h20763061C0630020806370760000098D81ADD00C5D8D31AC5D8C998CBECC5D8D;
defparam sp_inst_3.INIT_RAM_23 = 256'h2076306100003BFF4804040547FF4C04040553FF500404055FFF880404054076;
defparam sp_inst_3.INIT_RAM_24 = 256'h000000000000000000008400B2CCD98C008C9FFF807660767061806300204063;
defparam sp_inst_3.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_26 = 256'h0005759FB2CDFD8DB2CC00000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_27 = 256'h0000000000000000000000008400A2CCD98C008C6180008C57FF380467FF4804;
defparam sp_inst_3.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_29 = 256'h38040000759FA2CDFD8DA2CC0000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2A = 256'h000000000000000000000000000000000000840092CCD98C008CF59F008CA3FF;
defparam sp_inst_3.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2C = 256'h008CEBFF3C048C00040C759F92CDFD8D92CC0000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2D = 256'h00000000000000000000000000000000000000000000840082CCD98C008C6180;
defparam sp_inst_3.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2F = 256'hD98C008CF59F008C37FF3C040000759F82CDFD8D82CC00000000000000000000;
defparam sp_inst_3.INIT_RAM_30 = 256'h00000000000000000000000000000000000000000000000000000000840072CC;
defparam sp_inst_3.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_32 = 256'h840062CCD98C008C6180008C7FFF40042000140C759F72CDFD8D72CC00000000;
defparam sp_inst_3.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_35 = 256'h000000000000840052CCD98C008CF59F008CCBFF40040000759F62CDFD8D62CC;
defparam sp_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_37 = 256'h52CDFD8D52CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_38 = 256'h00000000000000000000840042CCD98C008C6180008C13FF4404B400240C759F;
defparam sp_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3A = 256'h0000759F42CDFD8D42CC00000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3B = 256'h00000000000000000000000000000000840032CCD98C008CF59F008C5FFF4404;
defparam sp_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3D = 256'h00053FFF4800340C759F32CDFD8D32CC00000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3E = 256'h000000000000000000000000840022CCD98C008C6180008C97FF3804A7FF4C04;
defparam sp_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_4 (
    .DO({sp_inst_4_dout_w[15:0],sp_inst_4_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_4}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_4.READ_MODE = 1'b0;
defparam sp_inst_4.WRITE_MODE = 2'b00;
defparam sp_inst_4.BIT_WIDTH = 16;
defparam sp_inst_4.BLK_SEL = 3'b001;
defparam sp_inst_4.RESET_MODE = "SYNC";
defparam sp_inst_4.INIT_RAM_00 = 256'h38040000759F22CDFD8D22CC0000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_01 = 256'h000000000000000000000000000000000000840012CCD98C008CF59F008CE3FF;
defparam sp_inst_4.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_03 = 256'h008C2BFF3C04CC00080C759F12CDFD8D12CC0000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_04 = 256'h00000000000000000000000000000000000000000000840002CCD98C008C6180;
defparam sp_inst_4.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_06 = 256'hD98C008CF59F008C77FF3C040000759F02CDFD8D02CC00000000000000000000;
defparam sp_inst_4.INIT_RAM_07 = 256'h000000000000000000000000000000000000000000000000000000008400F2CC;
defparam sp_inst_4.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_09 = 256'h8400E2CCD98C008C6180008CBFFF40046000180C759FF2CDFD8DF2CC00000000;
defparam sp_inst_4.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0C = 256'h0000000000008400D2CCD98C008CF59F008C0BFF40040000759FE2CDFD8DE2CC;
defparam sp_inst_4.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0E = 256'hD2CDFD8DD2CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0F = 256'h000000000000000000008400C2CCD98C008C6180008C53FF4404F400280C759F;
defparam sp_inst_4.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_11 = 256'h0000759FC2CDFD8DC2CC00000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_12 = 256'h000000000000000000000000000000008400B2CCD98C008CF59F008C9FFF4404;
defparam sp_inst_4.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_14 = 256'h00057FFF8800380C759FB2CDFD8DB2CC00000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_15 = 256'h0000000000000000000000008400A2CCD98C008C6180008CD7FF3804E7FF5004;
defparam sp_inst_4.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_17 = 256'h38040000759FA2CDFD8DA2CC0000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_18 = 256'h000000000000000000000000000000000000840092CCD98C008CF59F008C23FF;
defparam sp_inst_4.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1A = 256'h008C6BFF3C040C000C0C759F92CDFD8D92CC0000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1B = 256'h00000000000000000000000000000000000000000000840082CCD98C008C6180;
defparam sp_inst_4.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1D = 256'hD98C008CF59F008CB7FF3C040000759F82CDFD8D82CC00000000000000000000;
defparam sp_inst_4.INIT_RAM_1E = 256'h00000000000000000000000000000000000000000000000000000000840072CC;
defparam sp_inst_4.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_20 = 256'h840062CCD98C008C6180008CFFFF4004A0001C0C759F72CDFD8D72CC00000000;
defparam sp_inst_4.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_23 = 256'h000000000000840052CCD98C008CF59F008C4BFF40040000759F62CDFD8D62CC;
defparam sp_inst_4.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_25 = 256'h52CDFD8D52CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_26 = 256'h00000000000000000000840042CCD98C008C6180008C93FF440434002C0C759F;
defparam sp_inst_4.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_28 = 256'h0000759F42CDFD8D42CC00000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_29 = 256'h00000000000000000000000000000000840032CCD98C008CF59F008CDFFF4404;
defparam sp_inst_4.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_2B = 256'h0005BFFFC8003C0C759F32CDFD8D32CC00000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_2C = 256'h000000000000000000000000840022CCD98C008C6180008C17FF380427FF8804;
defparam sp_inst_4.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_2E = 256'h38040000759F22CDFD8D22CC0000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_2F = 256'h000000000000000000000000000000000000840012CCD98C008CF59F008C63FF;
defparam sp_inst_4.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_31 = 256'h008CABFF3C044C00100C759F12CDFD8D12CC0000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_32 = 256'h00000000000000000000000000000000000000000000840002CCD98C008C6180;
defparam sp_inst_4.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_34 = 256'hD98C008CF59F008CF7FF3C040000759F02CDFD8D02CC00000000000000000000;
defparam sp_inst_4.INIT_RAM_35 = 256'h000000000000000000000000000000000000000000000000000000008400F2CC;
defparam sp_inst_4.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_37 = 256'h8400E2CCD98C008C6180008C3FFF4004E000200C759FF2CDFD8DF2CC00000000;
defparam sp_inst_4.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_3A = 256'h0000000000008400D2CCD98C008CF59F008C8BFF40040000759FE2CDFD8DE2CC;
defparam sp_inst_4.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_3C = 256'hD2CDFD8DD2CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_3D = 256'h000000000000000000008400C2CCD98C008C6180008CD3FF44047400300C759F;
defparam sp_inst_4.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_3F = 256'h0000759FC2CDFD8DC2CC00000000000000000000000000000000000000000000;

SP sp_inst_5 (
    .DO({sp_inst_5_dout_w[15:0],sp_inst_5_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_5}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_5.READ_MODE = 1'b0;
defparam sp_inst_5.WRITE_MODE = 2'b00;
defparam sp_inst_5.BIT_WIDTH = 16;
defparam sp_inst_5.BLK_SEL = 3'b001;
defparam sp_inst_5.RESET_MODE = "SYNC";
defparam sp_inst_5.INIT_RAM_00 = 256'h000000000000000000000000000000008400B2CCD98C008CF59F008C1FFF4404;
defparam sp_inst_5.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_02 = 256'h0184000C0800400C759FB2CDFD8DB2CC00000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_03 = 256'h0020406320763061000043FF04040005407620763061C0630020806360767061;
defparam sp_inst_5.INIT_RAM_04 = 256'h80766076706180630020406320763061000013FF04040405407620763061C063;
defparam sp_inst_5.INIT_RAM_05 = 256'h0000000000000000000000000000000000008400B2CC958C016CE3FF8C040405;
defparam sp_inst_5.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_07 = 256'h958C016C37FF8C040005759FB2CDFD8DB2CC0000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_08 = 256'h000000000000000000000000000000000000000000000000000000008400A2CC;
defparam sp_inst_5.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_0A = 256'h000000000000840092CC958C016C8BFF8C040405759FA2CDFD8DA2CC00000000;
defparam sp_inst_5.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_0C = 256'h92CDFD8D92CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_0D = 256'hAFFF8C040405807660767061806300208063607670610000DFFF8C040005759F;
defparam sp_inst_5.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000008400B2CC798C088C;
defparam sp_inst_5.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_10 = 256'h0020806360767061000003FF8C040005759FB2CDFD8DB2CC0000000000000000;
defparam sp_inst_5.INIT_RAM_11 = 256'h0184B2CCB2C00800B2CC040C1180B1AC72CC018DDA0CB2C072C4C076B0764063;
defparam sp_inst_5.INIT_RAM_12 = 256'h018C0D8CD40C018D35CDB2CDDA0C018EDA0CB2C48076707680630020C063B076;
defparam sp_inst_5.INIT_RAM_13 = 256'hBECC008C80766076706180630020806370760000018D81AD05AD0D8CD40C818D;
defparam sp_inst_5.INIT_RAM_14 = 256'h93FF5004F7FF04048BFF47FF0184BECC9BFF57FF0004A7FF63FFE004E3FF0404;
defparam sp_inst_5.INIT_RAM_15 = 256'h3BFFF7FFE00477FF0404BECC008C807660767061806300208063607670610000;
defparam sp_inst_5.INIT_RAM_16 = 256'h0020806360767061000027FF50048BFF04041FFFDBFF0184BECC2FFFEBFF0004;
defparam sp_inst_5.INIT_RAM_17 = 256'h000000000000000000000000000000008400B2CC418C16CC8076607670618063;
defparam sp_inst_5.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_19 = 256'h6FFF800477FFB804759FB2CDFD8DB2CC00000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_1A = 256'h2FFFFC0437FF04043FFF000447FF40044FFF000457FF20045FFFC00467FF4004;
defparam sp_inst_5.INIT_RAM_1B = 256'hEFFF5404F7FF0004FFFF4C0407FF90040FFFFC0417FFA0041FFF980427FF8404;
defparam sp_inst_5.INIT_RAM_1C = 256'hAFFF3404B7FF8004BFFF6C04C7FF4804CFFF6804D7FF8804DFFF6404E7FFC004;
defparam sp_inst_5.INIT_RAM_1D = 256'hA2CCA2C5B2C48076607670618063002080636076706100009FFFBC04A7FF5004;
defparam sp_inst_5.INIT_RAM_1E = 256'h818CB2CC37FF0184818C418C818C3D8C818C918CB2CC5BFF0184818CC18C818C;
defparam sp_inst_5.INIT_RAM_1F = 256'h008CC076A076B06140630020806360767061000017FF0184818C058C818C398C;
defparam sp_inst_5.INIT_RAM_20 = 256'h7ECC1C00A2C0BBFF4004C3FF0004CBFF0184818CC18C818CB2CC6400B2C07ECC;
defparam sp_inst_5.INIT_RAM_21 = 256'hB0610000998D1C0CB2CDB2CC058CB2CCE18DFC0CA2CDA2CC058CA2CC13FF0184;
defparam sp_inst_5.INIT_RAM_22 = 256'hB0614063002040632076306100004FFF0004407620763061C0630020C063A076;
defparam sp_inst_5.INIT_RAM_23 = 256'hD800C58D080DB58D040D4ECCA2C0B2C092C04ECC00EC52C662C572C4C076A076;
defparam sp_inst_5.INIT_RAM_24 = 256'h2BFF72C462C562CC058C62CC72C0158DF80C72CD92CC818C018C31ACA2CC52CD;
defparam sp_inst_5.INIT_RAM_25 = 256'hB2CC058CB2CCE7FF0184018C31ACB2CC31AD31CC180C92CEF1AD00CD3C00B2C0;
defparam sp_inst_5.INIT_RAM_26 = 256'h52CD1C004D9F018C31ACA2CC52CDA2CC058CA2CC72CC198C72CCC18D140CB2CD;
defparam sp_inst_5.INIT_RAM_27 = 256'hB2C06FFF72C462C562CC058C62CC72C0158DE00C72CD92CC818C018C31ACA2CC;
defparam sp_inst_5.INIT_RAM_28 = 256'h1C0CB2CDB2CC058CB2CC2FFF0184018C31AC61AD00CD31ACB2CC918D92CC3800;
defparam sp_inst_5.INIT_RAM_29 = 256'h31ACE1AD00CD218C31ACB2CC918D92CC3C00B2C013FF72C40185058C62CCC58D;
defparam sp_inst_5.INIT_RAM_2A = 256'h52CDA2CC058CA2CC72CC218C72CCC18D1C0CB2CDB2CC058CB2CCCFFF0184018C;
defparam sp_inst_5.INIT_RAM_2B = 256'h62C572C4C076A076B06140630020C063A076B06100000000F19F018C31ACA2CC;
defparam sp_inst_5.INIT_RAM_2C = 256'h018C31ACA2CC11ADFF6D3800BEC047FF72C462C5A2CC958C5ECCBEC05ECC00CC;
defparam sp_inst_5.INIT_RAM_2D = 256'hEBFF72C40185058C62CCC58D3C0CBECDBECC058CBECCA2CC058CA2CC13FF0184;
defparam sp_inst_5.INIT_RAM_2E = 256'hBECDBECC058CBECCA2CC058CA2CCB7FF0184018C31ACA2CCA1ADFF6D3800BEC0;
defparam sp_inst_5.INIT_RAM_2F = 256'hB2C042C752C662C572C4C076A076B06140630020C063A076B0610000C58D3C0C;
defparam sp_inst_5.INIT_RAM_30 = 256'hB2CCB3FF01C462C50186818C31AC818C52CC818DB2CC31AE72CC918DB2CC4800;
defparam sp_inst_5.INIT_RAM_31 = 256'h62C572C40076E076F06100630020C063A076B0610000B5AC42CCB2CDB2CC058C;
defparam sp_inst_5.INIT_RAM_32 = 256'h62CC92CC058C8D8C42CC140092CC8D8C42CC15801D8C42CCB2C032C842C752C6;
defparam sp_inst_5.INIT_RAM_33 = 256'h5BFF0184018C31AC32CDB2CD058DB2CC3000A2CC72CC97FF72C492C5600092CC;
defparam sp_inst_5.INIT_RAM_34 = 256'h0063E076F06100009DAC42CC92CD92CC058C92CCCDAC52CCA2CDA2CC058CA2CC;
defparam sp_inst_5.INIT_RAM_35 = 256'h818C5ECCB2C0A2C05ACC01AC5ECC00ED00CC62C572C4C076A076B06140630020;
defparam sp_inst_5.INIT_RAM_36 = 256'h3800B2C0B3FF72C462C5BDAC400C5ACD62CC098C62CC72C0158DFC0C72CDA2CC;
defparam sp_inst_5.INIT_RAM_37 = 256'hC58D1C0CB2CDB2CC058CB2CC73FF0184018C31AC71AD00AD31ACB2CC918DA2CC;
defparam sp_inst_5.INIT_RAM_38 = 256'h018C31ACF1AD00AD218C31ACB2CC918DA2CC3C00B2C057FF72C40185058C62CC;
defparam sp_inst_5.INIT_RAM_39 = 256'h31AD00AD3C00B2C0FBFF72C462C55C00C18D1C0CB2CDB2CC058CB2CC13FF0184;
defparam sp_inst_5.INIT_RAM_3A = 256'h0000C18D140CB2CDB2CC058CB2CCB7FF0184018C31ACB2CC31AD31CC180CA2CE;
defparam sp_inst_5.INIT_RAM_3B = 256'hB2CC31AC72CCB2CD1400B2CC040C62C572C4C076B07640630020C063A076B061;
defparam sp_inst_5.INIT_RAM_3C = 256'h52C662C572C4C076A076B06140630020C063B0760184B2CCE59F62CDFD8D62CC;
defparam sp_inst_5.INIT_RAM_3D = 256'h008D5BFF28040185FD8C31ACB2CC4ECD0400B2C0A2C04ACC01AC4ECC010D00EC;
defparam sp_inst_5.INIT_RAM_3E = 256'h518DB2CC018DFD8C4ECC6580A2CC92CC000709A0B5CC280D000709A0358E52CC;
defparam sp_inst_5.INIT_RAM_3F = 256'h4BFF018462C5800601A74ACD31AC72CC31ADB2CC018D818C858C4ACC418092CC;

SP sp_inst_6 (
    .DO({sp_inst_6_dout_w[15:0],sp_inst_6_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_6}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_6.READ_MODE = 1'b0;
defparam sp_inst_6.WRITE_MODE = 2'b00;
defparam sp_inst_6.BIT_WIDTH = 16;
defparam sp_inst_6.BLK_SEL = 3'b001;
defparam sp_inst_6.RESET_MODE = "SYNC";
defparam sp_inst_6.INIT_RAM_00 = 256'h4ACE818CC18C818C92CC31AD72CC31ADB2CC018D818C858C4ACCA2CC040C5400;
defparam sp_inst_6.INIT_RAM_01 = 256'h0020C063A076B0610000F9ACB2CD4ECCB2CC058CB2CCF7FF01A462C5018601C7;
defparam sp_inst_6.INIT_RAM_02 = 256'h77FF4C04040583FF480404058FFF340404059BFF040404058076607670618063;
defparam sp_inst_6.INIT_RAM_03 = 256'h00053BFF9404040547FF9004040553FF8C0404055FFF880404056BFF50040405;
defparam sp_inst_6.INIT_RAM_04 = 256'h44040005FFFF400400050BFF3C04000517FF3804000523FF9C0404052FFF9804;
defparam sp_inst_6.INIT_RAM_05 = 256'h000000000000000000000000000000000000000000008400B2CCC98C0E2CF3FF;
defparam sp_inst_6.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_07 = 256'h040533FF940404053FFF90040405759FB2CDFD8DB2CC00000000000000000000;
defparam sp_inst_6.INIT_RAM_08 = 256'h70610000F7FF8C04000503FF9C0404050FFF980404051BFF3404040527FF0404;
defparam sp_inst_6.INIT_RAM_09 = 256'hB2CC958C016CDBFF018492CC9FFF018492CC8076607670618063002080636076;
defparam sp_inst_6.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000008400;
defparam sp_inst_6.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0C = 256'h016C07FF807660767061806300208063607670610000759FB2CDFD8DB2CC0000;
defparam sp_inst_6.INIT_RAM_0D = 256'h00000000000000000000000000000000000000000000000000008400B2CC958C;
defparam sp_inst_6.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0F = 256'h407620763061C06300208063607670610000759FB2CDFD8DB2CC000000000000;
defparam sp_inst_6.INIT_RAM_10 = 256'hF3FF1C005BFF93FFAFFF407620763061C0630020406320763061000043FF0804;
defparam sp_inst_6.INIT_RAM_11 = 256'h0000000000008400B2CC958C016C807660767061806300204063207630610000;
defparam sp_inst_6.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_13 = 256'hB2CDFD8DB2CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_14 = 256'h00000000000000000000000000000000000000008400A2CCED8C004CFC00759F;
defparam sp_inst_6.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_16 = 256'h0000840092CCED8C004C5800759FA2CDFD8DA2CC000000000000000000000000;
defparam sp_inst_6.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_18 = 256'h92CC000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_19 = 256'h00000000000000000000000000000000840082CCED8C004C2C00759F92CDFD8D;
defparam sp_inst_6.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_1B = 256'h6076706100008400759F82CDFD8D82CC00000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_1C = 256'h31AC000C5D8DF98C5D8C858C7ECCAEC07ECC008CC076A076B061406300208063;
defparam sp_inst_6.INIT_RAM_1D = 256'h818C058CCE0C0000F19F118C818C058CCE0C0000098DAACDCE0C83FFAACC5D8C;
defparam sp_inst_6.INIT_RAM_1E = 256'h058CCE0C0000F19F118C818C058CCE0C00000980CE0CAECC098CCE0CF19F058C;
defparam sp_inst_6.INIT_RAM_1F = 256'h0000000000000000000000008400B2CC080C4BFFAECC098CCE0CF19F058C818C;
defparam sp_inst_6.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_21 = 256'h0184AECC759FB2CDFD8DB2CC0000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_22 = 256'h818C858C7ECC7ACC01AC7ECC00AD008CC076A076B06140630020C063A076B061;
defparam sp_inst_6.INIT_RAM_23 = 256'h818C058CCE0C0000F19F118C818C058CCE0C0000098DAECDCE0C03FFAECCF98C;
defparam sp_inst_6.INIT_RAM_24 = 256'hCE0C0000F19F118C818C058CCE0C0000098D7ACDCE0CAACC098CCE0CF19F058C;
defparam sp_inst_6.INIT_RAM_25 = 256'h000000000000000000008400B2CC080CC7FFAACC098CCE0CF19F058C818C058C;
defparam sp_inst_6.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_27 = 256'h0000759FB2CDFD8DB2CC00000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_28 = 256'h01847ECCBEC07ACC01AC7ECC00AD008CC076A076B06140630020C063A076B061;
defparam sp_inst_6.INIT_RAM_29 = 256'hC063A076B061000027FF018401A57ECC818D5D8C31ACBECC7ACDBECC008CCBFF;
defparam sp_inst_6.INIT_RAM_2A = 256'hBECC008C57FF01847ECCBEC07ACC01AC7ECC00AD008CC076A076B06140630020;
defparam sp_inst_6.INIT_RAM_2B = 256'h0020C063A076B0610000ABFF018401A57ECC818D5D8CB1ACBECC5D8D300C7ACC;
defparam sp_inst_6.INIT_RAM_2C = 256'h0000000000000000000000008400B2CC880C13FF940404058076607670618063;
defparam sp_inst_6.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2E = 256'h94040005759FB2CDFD8DB2CC0000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000008400A2CC880C6BFF;
defparam sp_inst_6.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_31 = 256'h92CC880C1FFF04043C05C3FF94040405759FA2CDFD8DA2CC0000000000000000;
defparam sp_inst_6.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000008400;
defparam sp_inst_6.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_34 = 256'hA80434055FFFB00400056BFFB404780577FF4404F405759F92CDFD8D92CC0000;
defparam sp_inst_6.INIT_RAM_35 = 256'h60767061806300208063607670610184000C3BFF5404000547FFAC04F80553FF;
defparam sp_inst_6.INIT_RAM_36 = 256'h0000000000000000000000000000000000008400B2CC980C07FF540400058076;
defparam sp_inst_6.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_38 = 256'hAECCAECC008CDBFF5004759FB2CDFD8DB2CC0000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_39 = 256'h3061C06300208063607670610000AECC008CB3FF5404C3FF50040C0511800D8C;
defparam sp_inst_6.INIT_RAM_3A = 256'h008CC0769077A076B061406300204063207630610000F7FF50040C0540762076;
defparam sp_inst_6.INIT_RAM_3B = 256'h2D8D380D218D300D7ECCB6C0BAC0BECCF80C7ACC01AC7ECC42C852C700CD62C5;
defparam sp_inst_6.INIT_RAM_3C = 256'h0185818C31AC000CBACD00000800B6CCC00CBACCDC0C1C00B6CC400CBACC480C;
defparam sp_inst_6.INIT_RAM_3D = 256'h31AC62CDA2CC2C00A2C0ABFF2804000537FF0404000537FF100400054FFF0804;
defparam sp_inst_6.INIT_RAM_3E = 256'h300C7ECDDFFF040401857ECCD1ACA2CD7ACCA2CC058CA2CC07FF24040185018C;
defparam sp_inst_6.INIT_RAM_3F = 256'h2580A2CCA2CCFD8CA2CCB2CC008C2BFF1004A2CC018C026C47FF3404000511AC;

SP sp_inst_7 (
    .DO({sp_inst_7_dout_w[15:0],sp_inst_7_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_7}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_7.READ_MODE = 1'b0;
defparam sp_inst_7.WRITE_MODE = 2'b00;
defparam sp_inst_7.BIT_WIDTH = 16;
defparam sp_inst_7.BLK_SEL = 3'b001;
defparam sp_inst_7.RESET_MODE = "SYNC";
defparam sp_inst_7.INIT_RAM_00 = 256'h008CD3FF18041180A2CC5FFF34040005C19F818CB1ACB6CCB2CD1980058CB2CC;
defparam sp_inst_7.INIT_RAM_01 = 256'h8FFF2804CDAC300C7ECDBECCFC0C0D80058C818CB1ACBACCB2CDBEC0F5806D8C;
defparam sp_inst_7.INIT_RAM_02 = 256'h018D42CC31AD9ECC8D8DFD8CB2CC25809ECC9ECC1D8C008C7FFF3004B2CC008C;
defparam sp_inst_7.INIT_RAM_03 = 256'h2C00A2C0B2CC480C0D8D480CB2CDB2CC040C0D80B2CC018D42CC8D8DB2CC1400;
defparam sp_inst_7.INIT_RAM_04 = 256'hBECCF80C0C00D1ACA2CDB2CCA2CC058CA2CC02EC008CFBFF240431B752CDA2CC;
defparam sp_inst_7.INIT_RAM_05 = 256'hE076F06100630020C0639077A076B0610184BECC3FFF04040005CBFF30040005;
defparam sp_inst_7.INIT_RAM_06 = 256'hA2CE52CC3ECC63FF50040C05EFFF34041C05EFFF200420053ECC22C5008C0076;
defparam sp_inst_7.INIT_RAM_07 = 256'h52CD25AC400CA2CD3180BECCBECC008CCFFF30040185040601A701C852CC52CD;
defparam sp_inst_7.INIT_RAM_08 = 256'h006300200063E076F0610184BECCBECCF80C0C00018D56CD058C22CC018D22CC;
defparam sp_inst_7.INIT_RAM_09 = 256'h52CC4C0C13FF380400052BFF340400052BFF20042005B6C032C40076E076F061;
defparam sp_inst_7.INIT_RAM_0A = 256'hBAC08180BECCBECC008C03FF30040185080601A701C852CC52CDA2CE56CC800C;
defparam sp_inst_7.INIT_RAM_0B = 256'hB6CCB1ACB6CC918D31ACC2CDBACC018D91AD39ADC2CD31AC32CDBACCBACE4C00;
defparam sp_inst_7.INIT_RAM_0C = 256'h38040005BECCF80C0DACB6CD918C31ACC2CDBACCB18D0C0CBACDBACC058CBACC;
defparam sp_inst_7.INIT_RAM_0D = 256'hFBFF480450A5FF45BAC0807660767061806300200063E076F0610184BECCD3FF;
defparam sp_inst_7.INIT_RAM_0E = 256'h818D31AC280C818D818C918C018CD18CFF4C4980008CAFFF2084FF445D80008C;
defparam sp_inst_7.INIT_RAM_0F = 256'h7076806300208063607670610184BACCBACC31AC818C3D8C818C018C418CFF4C;
defparam sp_inst_7.INIT_RAM_10 = 256'h318DB2CC058D318CB2CC018DAECD358C31ADB2CD018CB2CCAECC00ACB2C48076;
defparam sp_inst_7.INIT_RAM_11 = 256'h118CB2CC418DB2CC418DB2CC058D418CB2CC3180B2CC0DAC118CB2CC318DB2CC;
defparam sp_inst_7.INIT_RAM_12 = 256'hB2CC0DAC118CB2CC218DB2CC218DB2CC058D218CB2CC418DB2CC118DB2CC458D;
defparam sp_inst_7.INIT_RAM_13 = 256'h63FF018401CC03FF63FF43FF9FFF807660767061806300208063707600002180;
defparam sp_inst_7.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000008400B2CCC98C0E2C;
defparam sp_inst_7.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_16 = 256'h0000000000008400A2CCC98C0E2C7FFF759FB2CDFD8DB2CC0000000000000000;
defparam sp_inst_7.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_18 = 256'hA2CDFD8DA2CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_19 = 256'h018DD58CFF2C018D008CA3FF6FFF0180498CFF2CADAC040C008DDBFF9804759F;
defparam sp_inst_7.INIT_RAM_1A = 256'h19AC040C018DB18CFF4C0180018C31ACA18C008C898DBDAC4C0D018C658CFF4C;
defparam sp_inst_7.INIT_RAM_1B = 256'h818CFF4C018D080DC58CFF4C29AC340C018D558CFF2C0180418CFF4C28000404;
defparam sp_inst_7.INIT_RAM_1C = 256'h018D200DA18CFF4C018D200DE58CFF4C39AC380C018D758CFF2C4C00018D080D;
defparam sp_inst_7.INIT_RAM_1D = 256'h29AC2C0C018DF58CFF2C0180E18CFF4C9000080419AC080C018D518CFF4C1400;
defparam sp_inst_7.INIT_RAM_1E = 256'h858CFF4C29AC300C018D158CFF2CBC00018D0C0D218CFF4C018D0C0D658CFF4C;
defparam sp_inst_7.INIT_RAM_1F = 256'h018D3C0DA58CFF4C29AC3C0C018D358CFF2C8400018D100D418CFF4C018D100D;
defparam sp_inst_7.INIT_RAM_20 = 256'h818CFF4C018D040DC58CFF4C39AC400C018D558CFF2C4C00018D3C0D618CFF4C;
defparam sp_inst_7.INIT_RAM_21 = 256'hC58CFF2C6C000180C18CFF4C8800100419AC0C0C018D318CFF4C1400018D040D;
defparam sp_inst_7.INIT_RAM_22 = 256'h100C018DA18CFF4CB800018D080DF18CFF4C018D080D358CFF4CDDAC400C018D;
defparam sp_inst_7.INIT_RAM_23 = 256'h018D080DA58CFF4C81AC400C018D358CFF2CAC000180318CFF4C2400140419AC;
defparam sp_inst_7.INIT_RAM_24 = 256'hFF2C0180A18CFF4CC0000C0419AC140C018D118CFF4C5C00018D080D618CFF4C;
defparam sp_inst_7.INIT_RAM_25 = 256'h018DD58CFF2C0400018D180DE18CFF4C018D180D258CFF4C29AC2C0C018DB58C;
defparam sp_inst_7.INIT_RAM_26 = 256'h29AC3C0C018DF58CFF2CCC00018D1C0D018CFF4C018D1C0D458CFF4C29AC300C;
defparam sp_inst_7.INIT_RAM_27 = 256'h858CFF4C81AC400C018D158CFF2C9400018D400D218CFF4C018D400D658CFF4C;
defparam sp_inst_7.INIT_RAM_28 = 256'h818CFF4CB800280419AC180C018DF18CFF4C5C00018D040D418CFF4C018D040D;
defparam sp_inst_7.INIT_RAM_29 = 256'hFF2C0400018D240DC18CFF4C018D240D058CFF4C29AC2C0C018D958CFF2C0180;
defparam sp_inst_7.INIT_RAM_2A = 256'h018DD58CFF2CCC00018D340DE18CFF4C018D340D258CFF4C29AC300C018DB58C;
defparam sp_inst_7.INIT_RAM_2B = 256'h81AC400C018DF58CFF2C9400018D140D018CFF4C018D140D458CFF4C29AC3C0C;
defparam sp_inst_7.INIT_RAM_2C = 256'hB0002C0419AC1C0C018DD18CFF4C5C00018D140D218CFF4C018D140D658CFF4C;
defparam sp_inst_7.INIT_RAM_2D = 256'h018D280DA18CFF4C018D280DE58CFF4C29AC2C0C018D758CFF2C0180618CFF4C;
defparam sp_inst_7.INIT_RAM_2E = 256'hFF0CCC00018D2C0DC18CFF4C018D2C0D058CFF4C29AC300C018D958CFF0C0400;
defparam sp_inst_7.INIT_RAM_2F = 256'h018DD58CFF0C9400018D140DE18CFF4C018D140D258CFF4C29AC3C0C018DB58C;
defparam sp_inst_7.INIT_RAM_30 = 256'h19AC200C018DB18CFF4C5C00018D140D018CFF4C018D140D458CFF4C81AC400C;
defparam sp_inst_7.INIT_RAM_31 = 256'hFF4C018D040DB58CFF4C25AC400C018D458CFF0CE4000180418CFF4CA8001C04;
defparam sp_inst_7.INIT_RAM_32 = 256'hFF0CE4000180B18CFF4C4400300419AC240C018D218CFF4C0000018D040D718C;
defparam sp_inst_7.INIT_RAM_33 = 256'h018D918CFF4CA400018D180DE18CFF4C018D180D258CFF4CC9AC400C018DB58C;
defparam sp_inst_7.INIT_RAM_34 = 256'h1C0D958CFF4C6DAC400C018D258CFF0C90000180218CFF4CE000340419AC280C;
defparam sp_inst_7.INIT_RAM_35 = 256'h0180918CFF4C7C00440419AC2C0C018D018CFF4C4800018D1C0D518CFF4C018D;
defparam sp_inst_7.INIT_RAM_36 = 256'hC58CFF0CF000018D300DD18CFF4C018D300D158CFF4C29AC340C018DA58CFF0C;
defparam sp_inst_7.INIT_RAM_37 = 256'h400C018DE58CFF0CB800018D1C0DF18CFF4C018D1C0D358CFF4C29AC380C018D;
defparam sp_inst_7.INIT_RAM_38 = 256'h38041DAC300C018DC18CFF4C8000018D1C0D118CFF4C018D1C0D558CFF4CA5AC;
defparam sp_inst_7.INIT_RAM_39 = 256'h818CFF4C018D1C0DC58CFF4C49AC400C018D558CFF0C0180418CFF4CAC00AC00;
defparam sp_inst_7.INIT_RAM_3A = 256'h018DD58CFF0C0180C18CFF4C4800400419AC340C018D318CFF4C2400018D1C0D;
defparam sp_inst_7.INIT_RAM_3B = 256'h29AC380C018DF58CFF0CCC00018D380D018CFF4C018D380D458CFF4C29AC340C;
defparam sp_inst_7.INIT_RAM_3C = 256'h858CFF4C81AC400C018D158CFF0C9400018D180D218CFF4C018D180D658CFF4C;
defparam sp_inst_7.INIT_RAM_3D = 256'hFF4C4800780038041DAC380C018DF18CFF4C5C00018D180D418CFF4C018D180D;
defparam sp_inst_7.INIT_RAM_3E = 256'h0000018D180DB18CFF4C018D180DF58CFF4C25AC400C018D858CFF0C0180718C;
defparam sp_inst_7.INIT_RAM_3F = 256'hFFFF018D040DB18CFF4C018D040DF58CFF4C140048042DAC3C0C018D618CFF4C;

SP sp_inst_8 (
    .DO({sp_inst_8_dout_w[15:0],sp_inst_8_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_8}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_8.READ_MODE = 1'b0;
defparam sp_inst_8.WRITE_MODE = 2'b00;
defparam sp_inst_8.BIT_WIDTH = 16;
defparam sp_inst_8.BLK_SEL = 3'b001;
defparam sp_inst_8.RESET_MODE = "SYNC";
defparam sp_inst_8.INIT_RAM_00 = 256'h818CFF4C9000018D080DD18CFF4C018D080D158CFF4CB5AC400C018DA58CFF0C;
defparam sp_inst_8.INIT_RAM_01 = 256'h440D958CFF4C29AC2C0C018D258CFF0C0180118CFF4C9C004C0419AC400C018D;
defparam sp_inst_8.INIT_RAM_02 = 256'hFF4C018D480DB58CFF4C29AC300C018D458CFF0C3800018D440D518CFF4C018D;
defparam sp_inst_8.INIT_RAM_03 = 256'h140D918CFF4C018D140DD58CFF4C29AC3C0C018D658CFF0C0000018D480D718C;
defparam sp_inst_8.INIT_RAM_04 = 256'h9000018D140DB18CFF4C018D140DF58CFF4CB5AC400C018D858CFF0CC800018D;
defparam sp_inst_8.INIT_RAM_05 = 256'h87FF018D400DB18CFF4C018D400DF58CFF4C940054042DAC440C018D618CFF4C;
defparam sp_inst_8.INIT_RAM_06 = 256'h818CFF4C2000018D400DD18CFF4C018D400D158CFF4C45AC400C018DA58CFF0C;
defparam sp_inst_8.INIT_RAM_07 = 256'h4C0D958CFF4C29AC340C018D258CFF0C0180118CFF4C1C00500419AC480C018D;
defparam sp_inst_8.INIT_RAM_08 = 256'hFF4C018D400DB58CFF4C29AC380C018D458CFF0CC800018D4C0D518CFF4C018D;
defparam sp_inst_8.INIT_RAM_09 = 256'h400D918CFF4C018D400DD58CFF4C7DAC400C018D658CFF0C9000018D400D718C;
defparam sp_inst_8.INIT_RAM_0A = 256'h818CFF2C018D400DC58CFF2C1BFF4C00380431AC4C0C018D418CFF4C5800018D;
defparam sp_inst_8.INIT_RAM_0B = 256'hE800018D400DB18CFF2C018D400DF58CFF2C0DAC400C018D858CFF0C018D400D;
defparam sp_inst_8.INIT_RAM_0C = 256'h818CFF2C018D040DC58CFF2CDFFF018D040D598CFF0C7FFF1980018CA98CFF0C;
defparam sp_inst_8.INIT_RAM_0D = 256'h0000CFFF0000D7FF0000DFFF0000E7FF0000EFFF0000F7FF0000FFFF018D040D;
defparam sp_inst_8.INIT_RAM_0E = 256'h00008FFF000097FF00009FFF0000A7FF0000AFFF0000B7FF0000BFFF0000C7FF;
defparam sp_inst_8.INIT_RAM_0F = 256'h008C80766076706180635FFF000067FF00006FFF000077FF00007FFF000087FF;
defparam sp_inst_8.INIT_RAM_10 = 256'h000540061407C108006867FF0180018C31AC418C006C898D7DAC540DBACCBACC;
defparam sp_inst_8.INIT_RAM_11 = 256'h1805380677FF78041805340687FF40041805200697FF000418051C0627FF7804;
defparam sp_inst_8.INIT_RAM_12 = 256'h0C0703FF58040805A0C6006608073FFF280400053C061C0703FF000067FFB804;
defparam sp_inst_8.INIT_RAM_13 = 256'h0807E7FFA004100524061007D7FF5804100500C60066080713FFA00408051806;
defparam sp_inst_8.INIT_RAM_14 = 256'h4C00A7FF200418052C060807BBFFA0041805E0060807ABFF5804180560C60066;
defparam sp_inst_8.INIT_RAM_15 = 256'h5804080580C60066080777FF18040005340608078BFF580400058C060C074FFF;
defparam sp_inst_8.INIT_RAM_16 = 256'hFFFF58041005A0C6006608073BFFE00408058C0608075BFFA004080518063BFF;
defparam sp_inst_8.INIT_RAM_17 = 256'hBFFF58041805B0C600660807FBFF200410058C0608070FFFA004100524060807;
defparam sp_inst_8.INIT_RAM_18 = 256'hAFFF28040005580663FF6000BBFF200418058C060807CFFFA0041805E0060807;
defparam sp_inst_8.INIT_RAM_19 = 256'h0C0067FF00041805B80608077BFFE804000518060C078FFF6804000584060807;
defparam sp_inst_8.INIT_RAM_1A = 256'h080538061007DFFFDC0037FF00041805B80608074BFF50040005580614070FFF;
defparam sp_inst_8.INIT_RAM_1B = 256'h8C060C07EBFF0004000558060C07AFFFAC0007FF3C040805740608071BFF3C04;
defparam sp_inst_8.INIT_RAM_1C = 256'h100757FF5400AFFF00041805B8060807C3FF8004000564060807D7FFC0040005;
defparam sp_inst_8.INIT_RAM_1D = 256'hA80610071BFF18007FFF7C04080580068FFF3C0408057C0693FF3C0408053806;
defparam sp_inst_8.INIT_RAM_1E = 256'h006608072BFFE00400058C0608074BFFA00400051806FFFFFC0057FF80040805;
defparam sp_inst_8.INIT_RAM_1F = 256'h70C600660807FBFF200408051806FFFFA0040805C0060807EFFF5804080550C6;
defparam sp_inst_8.INIT_RAM_20 = 256'hAFFF60041005C806BFFF200410051806C3FFA0041005CC060807B3FF58041005;
defparam sp_inst_8.INIT_RAM_21 = 256'h0005240608071FFF1C0077FFA00418059806080767FF5804180550C600660807;
defparam sp_inst_8.INIT_RAM_22 = 256'h0805C00608070BFF58040805C0C60066080747FF200400058C0608075BFFA004;
defparam sp_inst_8.INIT_RAM_23 = 256'h1005CC060807CBFF58041005D0C60066080707FF20040805640608071BFFA004;
defparam sp_inst_8.INIT_RAM_24 = 256'h58041805A0C600660807C3FFA0041005C806C7FF2004100564060807DBFFA004;
defparam sp_inst_8.INIT_RAM_25 = 256'h2004000518066FFFA0040005C006080733FF30008BFFA0041805980608077BFF;
defparam sp_inst_8.INIT_RAM_26 = 256'hD406D7FFD4002FFF100400056406080743FF90040005C006080707FF04006BFF;
defparam sp_inst_8.INIT_RAM_27 = 256'h7C06E7FF78040805C0060807ABFFA80003FFE0040805CC06080723FFA0040805;
defparam sp_inst_8.INIT_RAM_28 = 256'h00051806ABFF8C040005CC0608076FFF6C00D3FF380408058006E3FFF8040805;
defparam sp_inst_8.INIT_RAM_29 = 256'h13FF100077FFB0041805DC0687FF00041805D80697FF4C040005C806A7FF0C04;
defparam sp_inst_8.INIT_RAM_2A = 256'h1805D80637FF64040805C8063BFFE4040805640608074FFF64040805CC060807;
defparam sp_inst_8.INIT_RAM_2B = 256'h08056C060807EFFF64040805E0060807B3FFB00017FFB0041805DC0627FF0004;
defparam sp_inst_8.INIT_RAM_2C = 256'h00660807ABFF200400058C060807BFFFA0040005E006080783FF8000DBFFE404;
defparam sp_inst_8.INIT_RAM_2D = 256'h006608076BFF20040805E00608077FFFA0040805C00608076FFF5804080550C6;
defparam sp_inst_8.INIT_RAM_2E = 256'h1005C8062BFF20041005E00608073FFFA0041005CC0608072FFF5804100560C6;
defparam sp_inst_8.INIT_RAM_2F = 256'h080797FF9400EFFFA004180598060807DFFF5804180530C60066080727FFA004;
defparam sp_inst_8.INIT_RAM_30 = 256'h00041805D806BBFF64040805C806BFFFE4040805E0060807D3FF64040805CC06;
defparam sp_inst_8.INIT_RAM_31 = 256'h20040005E006080773FFA0040005C006080737FF34009BFFB0041805DC06ABFF;
defparam sp_inst_8.INIT_RAM_32 = 256'hF1808ACC8ACC008CB3FF80766076706180630020806360767061000000005FFF;
defparam sp_inst_8.INIT_RAM_33 = 256'h018D31CC898CB2CC71CEFF2E018D31AC898CC1ADFF2DFD8CB2CC4400B2CC100C;
defparam sp_inst_8.INIT_RAM_34 = 256'hEBFFB4040C050186140740088ACC018DB18CFF2C8ACDBC0CB2CCB2CCFD8CB2CC;
defparam sp_inst_8.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000008400A2CC918C1C6C;
defparam sp_inst_8.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_37 = 256'h0000840092CCD58C182C4BFF0BFF3C04759FA2CDFD8DA2CC0000000000000000;
defparam sp_inst_8.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_39 = 256'h92CC000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_3A = 256'h00208063607670610000018D180DF18CFF2C018D180D358CFF2C759F92CDFD8D;
defparam sp_inst_8.INIT_RAM_3B = 256'hB2CDB2CC058CB2CC018031AC898CB2CCB1ADFF2D2800B2C08076607670618063;
defparam sp_inst_8.INIT_RAM_3C = 256'h0000000000000000000000000000000000008400A2CCD58C182C2BFFD58D100C;
defparam sp_inst_8.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_3E = 256'hFF2C018D180DB58CFF2C759FA2CDFD8DA2CC0000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_3F = 256'h8ACC8ACC008C6FFFC076A076B061406300208063607670610000018D180D718C;

SP sp_inst_9 (
    .DO({sp_inst_9_dout_w[15:0],sp_inst_9_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_9}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_9.READ_MODE = 1'b0;
defparam sp_inst_9.WRITE_MODE = 2'b00;
defparam sp_inst_9.BIT_WIDTH = 16;
defparam sp_inst_9.BLK_SEL = 3'b001;
defparam sp_inst_9.RESET_MODE = "SYNC";
defparam sp_inst_9.INIT_RAM_00 = 256'hCBFFB7FF200489AC018C31CC898C72CCB1CEFF2E8ACD618D100C72CD72C07180;
defparam sp_inst_9.INIT_RAM_01 = 256'h000000000000000000000000000000000000000000008400B2CCE58C472C27FF;
defparam sp_inst_9.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_03 = 256'hA2CCE58C472CFFFF24044BFF83FF759FB2CDFD8DB2CC00000000000000000000;
defparam sp_inst_9.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000008400;
defparam sp_inst_9.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_06 = 256'h33FF1804BC00018D040DD58CFF2C018D040D118CFF2C759FA2CDFD8DA2CC0000;
defparam sp_inst_9.INIT_RAM_07 = 256'h00000000000000000000000000000000000000000000840092CC918C1C6C73FF;
defparam sp_inst_9.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_09 = 256'hC063A076B0610000000087FF1004759F92CDFD8D92CC00000000000000000000;
defparam sp_inst_9.INIT_RAM_0A = 256'hFF0C218D280C018D058CFEEC8180018C458CFEECA2C0C076A076B06140630020;
defparam sp_inst_9.INIT_RAM_0B = 256'h280C018DE58CFEEC018DD18CFF0C31AD280C018D218CFF0C818D0C0C018D318C;
defparam sp_inst_9.INIT_RAM_0C = 256'h058D018C618CFF0C018DD18CFF0C31AD018C118CFF0C018D81CC00070980B1AE;
defparam sp_inst_9.INIT_RAM_0D = 256'hB5CC280D92CE6400B2CCFD8C018CB18CFF0C92CC018C318CFF0C018D218CFF0C;
defparam sp_inst_9.INIT_RAM_0E = 256'h0C0542C604074008B58C8D8CB2CC92CC000709A035CC280D92CE42CC000709A0;
defparam sp_inst_9.INIT_RAM_0F = 256'h00000000000000000000840082CC298C02CC9D80B2CCB2CCFD8CB2CC63FF0184;
defparam sp_inst_9.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_11 = 256'hB2C0759F82CDFD8D82CC00000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_12 = 256'h058CB2CC07FF01840C05E0C600460807958C8D8C31ACB2CC018D118CFF0C4400;
defparam sp_inst_9.INIT_RAM_13 = 256'h818CFF0C018D31AC898CB2CC41ADFF0D4400B2C0B1AC018C018CFF0CB2CDB2CC;
defparam sp_inst_9.INIT_RAM_14 = 256'h79AC2C0C018DF58CFEECB98D100CB2CDB2CC058CB2CC1C00A2CC040C11AC018C;
defparam sp_inst_9.INIT_RAM_15 = 256'h000000000000000000000000840072CCE58C472C13FFB7FFA3FF2004A180A2CC;
defparam sp_inst_9.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_17 = 256'h37FF6FFF759F72CDFD8D72CC0000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000840062CCE58C472CEBFF2404;
defparam sp_inst_9.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1A = 256'h858CFF0C018D040DC18CFF0C759F62CDFD8D62CC000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1B = 256'h52CC918C1C6C43FF47FF07FF1804D4000180D18CFF0C0180418CFF0C018D040D;
defparam sp_inst_9.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000008400;
defparam sp_inst_9.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1E = 256'h018DD58CFEEC3FFF14040180A18CFF0C0180118CFF0C759F52CDFD8D52CC0000;
defparam sp_inst_9.INIT_RAM_1F = 256'hA0C600460807B58C8D8CB2CC3400B2C00180D18CFF0C0180418CFF0C61AC300C;
defparam sp_inst_9.INIT_RAM_20 = 256'hB06140630020C063A076B0610000C98D0C0CB2CDB2CC058CB2CCB3FF01840C05;
defparam sp_inst_9.INIT_RAM_21 = 256'h818D0C0C018D718CFEECCD8D280C018D458CFEEC4580018C858CFEECC076A076;
defparam sp_inst_9.INIT_RAM_22 = 256'h81CC00070980B1AE280C018D258CFEEC018D118CFEEC31AD280C018D618CFEEC;
defparam sp_inst_9.INIT_RAM_23 = 256'hFEEC018D618CFEEC058D018CA18CFEEC018D118CFEEC31AD018C518CFEEC018D;
defparam sp_inst_9.INIT_RAM_24 = 256'hA2CE6ECC000709A0B5CC280DA2CE6C00B2CCFD8C018CF18CFEECA2CC018C718C;
defparam sp_inst_9.INIT_RAM_25 = 256'hABFF01A40C050186040740086ECC018DB58C8D8CB2CCA2CC000709A035CC280D;
defparam sp_inst_9.INIT_RAM_26 = 256'h0000000000000000000000000000840092CC518C05AC9580B2CCB2CCFD8CB2CC;
defparam sp_inst_9.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_28 = 256'h018DD58CFEEC759F92CDFD8D92CC000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_29 = 256'h140D918CFF0C018D140DD58CFF0C8FFF2004E9AC5C0C018D418CFEECE5AC2C0C;
defparam sp_inst_9.INIT_RAM_2A = 256'h00000000000000000000000000000000000000000000840082CC918C1C6C018D;
defparam sp_inst_9.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2C = 256'hEC000180618CFEEC0180D18CFEEC759F82CDFD8D82CC00000000000000000000;
defparam sp_inst_9.INIT_RAM_2D = 256'h00000000000000000000000000000000840072CC918C1C6CE7FFA7FF18044FFF;
defparam sp_inst_9.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2F = 256'h018D200DA58CFF0C759F72CDFD8D72CC00000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_30 = 256'hFEEC61AC300C018D058CFECC0180B18CFEEC0180218CFEEC018D200D618CFF0C;
defparam sp_inst_9.INIT_RAM_31 = 256'h3FFF01840C05D0C600460807B58C8D8CB2CC3400B2C00180018CFEEC0180718C;
defparam sp_inst_9.INIT_RAM_32 = 256'hFECC80766076706180630020C063A076B0610000C98D0C0CB2CDB2CC058CB2CC;
defparam sp_inst_9.INIT_RAM_33 = 256'h018D918CFEEC818D0C0C018DA18CFEEC2D8D280C018D758CFECC1580018CB58C;
defparam sp_inst_9.INIT_RAM_34 = 256'h818CFEEC018D81CC00070980B1AE280C018D558CFECC018D418CFEEC31AD280C;
defparam sp_inst_9.INIT_RAM_35 = 256'hA2CC018CA18CFEEC018D918CFEEC058D018CD18CFEEC018D418CFEEC31AD018C;
defparam sp_inst_9.INIT_RAM_36 = 256'h09A035CC280DA2CE8ECC000709A0B5CC280DA2CE6C00B2CCFD8C018C218CFEEC;
defparam sp_inst_9.INIT_RAM_37 = 256'hB2CCFD8CB2CC37FF01A40C050186040740088ECC018DB58C8D8CB2CCA2CC0007;
defparam sp_inst_9.INIT_RAM_38 = 256'h31AC898C01ADFF0DFD8CB2CC4400B2CC100C55AC2C0C018D858CFECC9580B2CC;
defparam sp_inst_9.INIT_RAM_39 = 256'hFF0C018DA18CFEECBC0CB2CCB2CCFD8CB2CC018D31CC898CB2CCB1CEFF0E018D;
defparam sp_inst_9.INIT_RAM_3A = 256'h0000840092CC918C1C6C47FF3C0493FF0180D18CFEEC0180418CFEEC018DD18C;
defparam sp_inst_9.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3C = 256'h92CC000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3D = 256'h61AC300C018DF58CFECC018D1C0DF18CFF0C018D1C0D358CFF0C759F92CDFD8D;
defparam sp_inst_9.INIT_RAM_3E = 256'h01840C05C0C600460807B58C8D8CB2CC3400B2C00180F18CFEEC0180618CFEEC;
defparam sp_inst_9.INIT_RAM_3F = 256'hB2C080767076806300208063607670610000C98D0C0CB2CDB2CC058CB2CCFBFF;

SP sp_inst_10 (
    .DO({sp_inst_10_dout_w[15:0],sp_inst_10_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_10}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_10.READ_MODE = 1'b0;
defparam sp_inst_10.WRITE_MODE = 2'b00;
defparam sp_inst_10.BIT_WIDTH = 16;
defparam sp_inst_10.BLK_SEL = 3'b001;
defparam sp_inst_10.RESET_MODE = "SYNC";
defparam sp_inst_10.INIT_RAM_00 = 256'hA2CC918C1C6CD58D100CB2CDB2CC058CB2CC018031AC898CB2CCB1ADFF0D2800;
defparam sp_inst_10.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000008400;
defparam sp_inst_10.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_03 = 256'h806370760000018D1C0DD18CFF0C018D1C0D158CFF0C759FA2CDFD8DA2CC0000;
defparam sp_inst_10.INIT_RAM_04 = 256'h000037FF8184D60C04058FFF708400445005A0C60046407620763061C0630020;
defparam sp_inst_10.INIT_RAM_05 = 256'hD60C080543FF408400446405D0C60046407620763061C0630020406320763061;
defparam sp_inst_10.INIT_RAM_06 = 256'h10840044780500C60046407620763061C06300204063207630610000EBFF8184;
defparam sp_inst_10.INIT_RAM_07 = 256'h30C60046407620763061C063002040632076306100009FFF8184D60C1005F7FF;
defparam sp_inst_10.INIT_RAM_08 = 256'h20763061C0630020406320763061000053FF8184D60C2005ABFFE08400448C05;
defparam sp_inst_10.INIT_RAM_09 = 256'h0020406320763061000007FF8184D60C40055FFFB0840044A00560C600464076;
defparam sp_inst_10.INIT_RAM_0A = 256'h30610000BBFF8184D60C800513FF80840044B40590C60046407620763061C063;
defparam sp_inst_10.INIT_RAM_0B = 256'h8184D60C0005C7FF50840044C805C0C60046407620763061C063002040632076;
defparam sp_inst_10.INIT_RAM_0C = 256'h7BFF20840044E005F0C60046407620763061C063002040632076306100006FFF;
defparam sp_inst_10.INIT_RAM_0D = 256'hF40520C60046407620763061C0630020406320763061000023FF8184D60C0005;
defparam sp_inst_10.INIT_RAM_0E = 256'h407620763061C06300204063207630610000D7FF8184D60C00052FFFF0840044;
defparam sp_inst_10.INIT_RAM_0F = 256'hC063002040632076306100008BFF8184D60C0005E3FFC08400240C0550C60046;
defparam sp_inst_10.INIT_RAM_10 = 256'h2076306100003FFF8184D60C000597FF90840024240580C60046407620763061;
defparam sp_inst_10.INIT_RAM_11 = 256'hF3FF8184D60C00054BFF608400243C05B0C60046407620763061C06300204063;
defparam sp_inst_10.INIT_RAM_12 = 256'h0025FFFF308400245005E0C60046407620763061C06300204063207630610000;
defparam sp_inst_10.INIT_RAM_13 = 256'h0024640510C60046407620763061C06300204063207630610000A7FF8184D60C;
defparam sp_inst_10.INIT_RAM_14 = 256'h0046407620763061C063002040632076306100005BFF8184D60C0045B3FF0084;
defparam sp_inst_10.INIT_RAM_15 = 256'h3061C063002040632076306100000FFF8184D60C008567FFD08400247C0540C6;
defparam sp_inst_10.INIT_RAM_16 = 256'h4063207630610000C3FF8184D60C01051BFFA0840024940570C6004640762076;
defparam sp_inst_10.INIT_RAM_17 = 256'h000077FF8184D60C0205CFFF70840024B005A0C60046407620763061C0630020;
defparam sp_inst_10.INIT_RAM_18 = 256'hD60C040583FF40840024C805D0C60046407620763061C0630020406320763061;
defparam sp_inst_10.INIT_RAM_19 = 256'h10840024E00500C60046407620763061C063002040632076306100002BFF8184;
defparam sp_inst_10.INIT_RAM_1A = 256'h30C60046407620763061C06300204063207630610000DFFF8184D60C080537FF;
defparam sp_inst_10.INIT_RAM_1B = 256'h20763061C0630020406320763061000093FF8184D60C1005EBFFE0840024F805;
defparam sp_inst_10.INIT_RAM_1C = 256'h0020406320763061000047FF8184D60C20059FFFB0840024100560C600464076;
defparam sp_inst_10.INIT_RAM_1D = 256'h30610000FBFF8184D60C400553FF80840024240590C60046407620763061C063;
defparam sp_inst_10.INIT_RAM_1E = 256'h8184D60C800507FF508400243805C0C60026407620763061C063002040632076;
defparam sp_inst_10.INIT_RAM_1F = 256'hBBFF208400245005F0C60026407620763061C06300204063207630610000AFFF;
defparam sp_inst_10.INIT_RAM_20 = 256'h680520C60026407620763061C0630020406320763061000063FF8184D60C0005;
defparam sp_inst_10.INIT_RAM_21 = 256'h407620763061C0630020406320763061000017FF8184D60C00056FFFF0840024;
defparam sp_inst_10.INIT_RAM_22 = 256'hC06300204063207630610000CBFF8184D60C000523FFC0840024800550C60026;
defparam sp_inst_10.INIT_RAM_23 = 256'h2076306100007FFF8184D60C0005D7FF90840024980580C60026407620763061;
defparam sp_inst_10.INIT_RAM_24 = 256'h33FF8184D60C00058BFF60840024B005B0C60026407620763061C06300204063;
defparam sp_inst_10.INIT_RAM_25 = 256'h00053FFF30840024C805E0C60026407620763061C06300204063207630610000;
defparam sp_inst_10.INIT_RAM_26 = 256'h0024E40510C60026407620763061C06300204063207630610000E7FF8184D60C;
defparam sp_inst_10.INIT_RAM_27 = 256'h0026407620763061C063002040632076306100009BFF8184D60C0005F3FF0084;
defparam sp_inst_10.INIT_RAM_28 = 256'h3061C063002040632076306100004FFF8184D60C0005A7FFD0840024FC0540C6;
defparam sp_inst_10.INIT_RAM_29 = 256'h406320763061000003FF8184D60C00055BFFA0840024140570C6002640762076;
defparam sp_inst_10.INIT_RAM_2A = 256'hD60CFFFF30840024C40560C60026018D000DF18CD60C80766076706180630020;
defparam sp_inst_10.INIT_RAM_2B = 256'hB2CCA2CD4000B2C00000A2CCB1AC92CCA2CD92CC018C818CD60CA2CC318C818C;
defparam sp_inst_10.INIT_RAM_2C = 256'hBD8D7C0CB2CDB2CC058CB2CC0181018C31AC898CB2CCB1AD002D2180058CB1AC;
defparam sp_inst_10.INIT_RAM_2D = 256'h018C118CD60C018D020DF18CD60C807660767061806300208063607670610000;
defparam sp_inst_10.INIT_RAM_2E = 256'h818CC18C018C118CD68C80766076706180630020806360767061000083FFB2CC;
defparam sp_inst_10.INIT_RAM_2F = 256'h018D3C0D118CD68C018D040DF18CD60CB6CC3D8C818C018C118CD68CBACCFD8C;
defparam sp_inst_10.INIT_RAM_30 = 256'h080DF18CD60C80767076806300208063607670610000A7FFF08400240185BACC;
defparam sp_inst_10.INIT_RAM_31 = 256'h018C118CD60C80766076706180630020806370760000BECC018C098CD18C018D;
defparam sp_inst_10.INIT_RAM_32 = 256'h898DB2CC718D400CB2CD018DB5CDF00DF18CD60C018E118CD60CB2CC7D8CCD8C;
defparam sp_inst_10.INIT_RAM_33 = 256'hD60CBFFF708400243C000180118CD60CDBFF408400240180018C31ACE18C002C;
defparam sp_inst_10.INIT_RAM_34 = 256'h80630020806360767061000000000800018DB5CDFDADFEED118CD60C018E118C;
defparam sp_inst_10.INIT_RAM_35 = 256'h13FF00041980008CD7FF00042980058CBECCBECC018C158CD40C807660767061;
defparam sp_inst_10.INIT_RAM_36 = 256'h018D100D0D8CD40CCBFF0184BACCBACC018CD10C2D80118CBECC2FFFC0840024;
defparam sp_inst_10.INIT_RAM_37 = 256'hFC0D0D8CD40C018D200D0D8CD40C97FF0184B6CCB6CC018CD00C2D80218CBECC;
defparam sp_inst_10.INIT_RAM_38 = 256'h0000F3FF83FFB084002423FF407620763061C06300208063607670610000018D;
defparam sp_inst_10.INIT_RAM_39 = 256'h15EC16F016F016F016F016F016F016F016F016F016F015D40020406320763061;
defparam sp_inst_10.INIT_RAM_3A = 256'h16F016F016F016F016F016F016F0167416741674167416741674167416741674;
defparam sp_inst_10.INIT_RAM_3B = 256'h16F016F016F016F016F016F016F016F016F016F016F016F016F016F016F016F0;
defparam sp_inst_10.INIT_RAM_3C = 256'h16F016F016F016F016F016F016F016F016F016F016F016F016F016F016F016F0;
defparam sp_inst_10.INIT_RAM_3D = 256'h159C152C16F016F016F016F016F016F016F016F016F016F014F4148C156416F0;
defparam sp_inst_10.INIT_RAM_3E = 256'hCAD3B0DDCA2000002020204B20202020159C16F016F014BC16F0146016F016F0;
defparam sp_inst_10.INIT_RAM_3F = 256'hB5ABBBC9CCC6D6200000A7CABCCDB8D6BCC20000D6CABBC3F7C6ABB40000CEED;

SP sp_inst_11 (
    .DO({sp_inst_11_dout_w[15:0],sp_inst_11_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_11}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_11.READ_MODE = 1'b0;
defparam sp_inst_11.WRITE_MODE = 2'b00;
defparam sp_inst_11.BIT_WIDTH = 16;
defparam sp_inst_11.BLK_SEL = 3'b001;
defparam sp_inst_11.RESET_MODE = "SYNC";
defparam sp_inst_11.INIT_RAM_00 = 256'h0000C9ABB5F7CCC6D6200000D2C2F1CFC6CE20200000BAABBBAACCC6D6200000;
defparam sp_inst_11.INIT_RAM_01 = 256'hD8B50000B0A7B2CFD5D820200000CEB8B5F7CBD0C32000002020A5C6C6CE2020;
defparam sp_inst_11.INIT_RAM_02 = 256'hF8C7BABB0000B0A7BFC6D6D5C7200000DCB0E5B0FDB320200000B6B7ACB3F2D0;
defparam sp_inst_11.INIT_RAM_03 = 256'hE6B4A7D02020000020F3B4E5B6B420200000EDB4485346B4B6200000A7D0DECE;
defparam sp_inst_11.INIT_RAM_04 = 256'h2020E2BFB8D620200000CEEDC2B3B1C2BC200000CEEDC8DAC6E6BC200000C5BA;
defparam sp_inst_11.INIT_RAM_05 = 256'h2F902EA82DE82D3C44490000CED0C2CFC8D8B72000002020EDB4D8B520200000;
defparam sp_inst_11.INIT_RAM_06 = 256'h2241004100000305502236000864122A2400147F000700002F00000000003064;
defparam sp_inst_11.INIT_RAM_07 = 256'h18004541464942007F423E453E000810000000000808006000003E0814081400;
defparam sp_inst_11.INIT_RAM_08 = 256'h08140000141400410800365600000000494936493600097130493C004545107F;
defparam sp_inst_11.INIT_RAM_09 = 256'h7F417F087F00494101097F0049491C227F00414136497F0011123E5132005101;
defparam sp_inst_11.INIT_RAM_0A = 256'h0100494946297F00514106097F0041417F107F000C0240407F001408013F2000;
defparam sp_inst_11.INIT_RAM_0B = 256'h040204004141552A5500417F4345610070086314630038401F201F0040400101;
defparam sp_inst_11.INIT_RAM_0C = 256'h7D4478047F00A4A40201080054547F483800444438447F005454000400004040;
defparam sp_inst_11.INIT_RAM_0D = 256'h0400545408047C0024241824FC00444478047C001804004000002810007D4000;
defparam sp_inst_11.INIT_RAM_0E = 256'h000000000000000000001414444C4400A0A04428440030401C201C0040402040;
defparam sp_inst_11.INIT_RAM_0F = 256'h08F01E21180030087000043F3F0478C0C040000000000C101000003000000000;
defparam sp_inst_11.INIT_RAM_10 = 256'h0200201800000418000000000000000016102719211E0070F000211E210018E0;
defparam sp_inst_11.INIT_RAM_11 = 256'h00000000B08000000000010101010000000002010202408040400007400000E0;
defparam sp_inst_11.INIT_RAM_12 = 256'h100010200F001008E00000016000608000000000300000000000010101000000;
defparam sp_inst_11.INIT_RAM_13 = 256'hF8003F240700F810000011201800488830002122300088087000202020000000;
defparam sp_inst_11.INIT_RAM_14 = 256'hE00022211C00880870000000000038C8380011200F001888E000112019000888;
defparam sp_inst_11.INIT_RAM_15 = 256'h4040100801001020000000000000000000000030000000C00000112200001008;
defparam sp_inst_11.INIT_RAM_16 = 256'h00001423180710E830C001360000080870000204200080400800040404044040;
defparam sp_inst_11.INIT_RAM_17 = 256'hF80810203F201008F80810201807080830C011203F207088F80827023C2000E0;
defparam sp_inst_11.INIT_RAM_18 = 256'h080021013F200800F8081E221807380830C000033F2008E8F80820233F2008E8;
defparam sp_inst_11.INIT_RAM_19 = 256'hF80820203F200000F80838263F201828F808007F80C008F80000202020000808;
defparam sp_inst_11.INIT_RAM_1A = 256'h10E001013F200808F8081020100F100810E018073F200800F8083F003F20F8F8;
defparam sp_inst_11.INIT_RAM_1B = 256'hF808002000000808081822213800080870000C033F208888F8085038180F1008;
defparam sp_inst_11.INIT_RAM_1C = 256'h38082C033020688018083C073C03080008F8010E0000C800780820201F000800;
defparam sp_inst_11.INIT_RAM_1D = 256'h02003806000000000C0040400000020200002020382038C808100020000038C8;
defparam sp_inst_11.INIT_RAM_1E = 256'h0000000000000000020080808080000000000000000002020000007F400000FE;
defparam sp_inst_11.INIT_RAM_1F = 256'h000010200E008880000020200E008080000011203F000080F808222219008080;
defparam sp_inst_11.INIT_RAM_20 = 256'h800020003F208080F80893946B0080800000202020008888800022221F008080;
defparam sp_inst_11.INIT_RAM_21 = 256'h80802020200000000800302D3F208080F8087F80C00098980000202020000000;
defparam sp_inst_11.INIT_RAM_22 = 256'h00001120FF800080808020201F008080000020003F2080808080203F3F208080;
defparam sp_inst_11.INIT_RAM_23 = 256'h8080202000008080800024243300808000000020202080808080A0200E008080;
defparam sp_inst_11.INIT_RAM_24 = 256'h8080310E200080808000300C300F80008080060801008000808010201F008000;
defparam sp_inst_11.INIT_RAM_25 = 256'h020000FF000000FF00003F0000007C8000002122210080808000061881808000;
defparam sp_inst_11.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000002020600000040000080;
defparam sp_inst_11.INIT_RAM_27 = 256'h0000000000000080C0C080800000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_28 = 256'h000000000000000000000000F0FE03010101FFFC000000000000000000000000;
defparam sp_inst_11.INIT_RAM_29 = 256'h7F7F07000000000000000000000000000000FEFFFFFF0F0FFFFFFFFF00000000;
defparam sp_inst_11.INIT_RAM_2A = 256'h00000000000000000000000000000000000000000000000000003F7FFFFFFFFF;
defparam sp_inst_11.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2C = 256'h7FC07F5C7E8C7E287D587CF47C907C2C7B247A1C791478B0784C774476AC834C;
defparam sp_inst_11.INIT_RAM_2D = 256'h86B08680862C8540848C84288C880020002A2E332E322E31828881B881408038;
defparam sp_inst_11.INIT_RAM_2E = 256'h0A0D8C588BF88B0C8ADC8A7C8A2089E489B88988895C887087908774873886E0;
defparam sp_inst_11.INIT_RAM_2F = 256'h2E2E2E2E2E2E544E54462E2E2E2E2E2E2E0A00003E2073256E756425656E2020;
defparam sp_inst_11.INIT_RAM_30 = 256'h2E2E4C495F542E2E2E2E2E2E2E0A000A7830656E68434B3A49686F742D0A0D0A;
defparam sp_inst_11.INIT_RAM_31 = 256'h69546C6168706550000D2E2E2E2E2E2E2E432E2E2E2E2E2E2E0A0D0A2E2E2E2E;
defparam sp_inst_11.INIT_RAM_32 = 256'hA150A104000A747072656920656C726554206F4300002E7472726E6961652072;
defparam sp_inst_11.INIT_RAM_33 = 256'hA610A5C4A578A52CA4E0A494A448A3FCA3B0A364A318A2CCA280A234A1E8A19C;
defparam sp_inst_11.INIT_RAM_34 = 256'hACD4AD24AA38A9ECA9A0A954A908A8BCA870A824A7D8A78CA740A6F4A6A8A65C;
defparam sp_inst_11.INIT_RAM_35 = 256'h7865ACF0AD24AD24AD24AD24AD24AD24AD24AD24AD24AD24AD24AD24AD24AD24;
defparam sp_inst_11.INIT_RAM_36 = 256'h61687269616F675F7865656C61687269616F675F7865656C61687269616F675F;
defparam sp_inst_11.INIT_RAM_37 = 256'h616F675F7865656C61687269616F675F7865656C61687269616F675F7865656C;
defparam sp_inst_11.INIT_RAM_38 = 256'h7865656C61687269616F675F7865656C61687269616F675F7865656C61687269;
defparam sp_inst_11.INIT_RAM_39 = 256'h61687269626F675F7865656C61687269626F675F7865656C61687269626F675F;
defparam sp_inst_11.INIT_RAM_3A = 256'h626F675F7865656C61687269626F675F7865656C61687269626F675F7865656C;
defparam sp_inst_11.INIT_RAM_3B = 256'h7865656C61687269626F675F7865656C61687269626F675F7865656C61687269;
defparam sp_inst_11.INIT_RAM_3C = 256'h61687269636F675F7865656C61687269636F675F7865656C61687269636F675F;
defparam sp_inst_11.INIT_RAM_3D = 256'h636F675F7865656C61687269636F675F7865656C61687269636F675F7865656C;
defparam sp_inst_11.INIT_RAM_3E = 256'h7865656C61687269636F675F7865656C61687269636F675F7865656C61687269;
defparam sp_inst_11.INIT_RAM_3F = 256'h61687269646F675F7865656C61687269646F675F7865656C61687269646F675F;

SP sp_inst_12 (
    .DO({sp_inst_12_dout_w[15:0],sp_inst_12_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_12}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_12.READ_MODE = 1'b0;
defparam sp_inst_12.WRITE_MODE = 2'b00;
defparam sp_inst_12.BIT_WIDTH = 16;
defparam sp_inst_12.BLK_SEL = 3'b001;
defparam sp_inst_12.RESET_MODE = "SYNC";
defparam sp_inst_12.INIT_RAM_00 = 256'h646F675F7865656C61687269646F675F7865656C61687269646F675F7865656C;
defparam sp_inst_12.INIT_RAM_01 = 256'h7865656C61687269646F675F7865656C61687269646F675F7865656C61687269;
defparam sp_inst_12.INIT_RAM_02 = 256'h321E941048001B0000000001FFFF035003680344000C034C032C0000656C6168;
defparam sp_inst_12.INIT_RAM_03 = 256'h0000F80082847E009252FF0082847F004A48CC0800004949494900007E427E00;
defparam sp_inst_12.INIT_RAM_04 = 256'hA62A0000884909094909880844241424147F44407F8000000000FF00FE020202;
defparam sp_inst_12.INIT_RAM_05 = 256'h404040404040000F80126722C8A899A80030302046230202420B420000011121;
defparam sp_inst_12.INIT_RAM_06 = 256'h242410200909090A893F60801E2292222CF41020001002000000000040444444;
defparam sp_inst_12.INIT_RAM_07 = 256'hC444840400F84242434102029444244404E48C104F20102011210101E628202C;
defparam sp_inst_12.INIT_RAM_08 = 256'h242410200909090A893F60801E2292222CF41020408808083F10010280FE82F2;
defparam sp_inst_12.INIT_RAM_09 = 256'h575517008041102C8890000020A08282400040404F20102011210101E628202C;
defparam sp_inst_12.INIT_RAM_0A = 256'h50004040007F15150010000044547F5444004240404055555555404017155755;
defparam sp_inst_12.INIT_RAM_0B = 256'h2CF410201012FF12100082428086A252820010105C5040405020400040487F48;
defparam sp_inst_12.INIT_RAM_0C = 256'hF80808084F20102011210101E628202C242410200909090A893F60801E229222;
defparam sp_inst_12.INIT_RAM_0D = 256'h4400424040200300103F20001611FF1090901010000080400718800008088888;
defparam sp_inst_12.INIT_RAM_0E = 256'h010000007F80FF9200051909D008D15210086888007F15150010000044547F54;
defparam sp_inst_12.INIT_RAM_0F = 256'hC444840400F84242434102029444244404E48C1080400300030C4080000000E0;
defparam sp_inst_12.INIT_RAM_10 = 256'h242410200909090A893F60801E2292222CF41020408808083F10010280FE82F2;
defparam sp_inst_12.INIT_RAM_11 = 256'hFE02FE0081410D030D11818100101010101040004F20102011210101E628202C;
defparam sp_inst_12.INIT_RAM_12 = 256'h080808084126214020106080C80AFF0888880000402116216710478010F017D8;
defparam sp_inst_12.INIT_RAM_13 = 256'h2222000081812F1181800000E424FF24E40460803F40010E88083010F010FF10;
defparam sp_inst_12.INIT_RAM_14 = 256'h8484840400004A4A4A4A0000A22AA3A4AAA66488007F02020202608000FE2222;
defparam sp_inst_12.INIT_RAM_15 = 256'h00004040804F10102040808000C05252525200004444444410106020FE929292;
defparam sp_inst_12.INIT_RAM_16 = 256'h00004040FC40404040407C0000FC4040404000005845404440204000807FC949;
defparam sp_inst_12.INIT_RAM_17 = 256'h9C642404007F27242720000000FEF212F2020000504845485820400062A324A4;
defparam sp_inst_12.INIT_RAM_18 = 256'hC05840404344404240204000FC04000200004040402001064C8208101828C80F;
defparam sp_inst_12.INIT_RAM_19 = 256'h000040407F21212100FF1F000808180F40FFF80040403F00071880804046C040;
defparam sp_inst_12.INIT_RAM_1A = 256'h10006010007F27242720000000FEF212F2020000504845485820400062A324A4;
defparam sp_inst_12.INIT_RAM_1B = 256'hA42400007F207F0080404080F808F8001010101009047F802100040412921E32;
defparam sp_inst_12.INIT_RAM_1C = 256'h2086FE00007F15150000040444547F5444006010101212FF12133040242424A6;
defparam sp_inst_12.INIT_RAM_1D = 256'h494900007840404040400000000082828282000031097F811127FF002010E324;
defparam sp_inst_12.INIT_RAM_1E = 256'h9010101000004444444401018242220622420200818989894121418100004949;
defparam sp_inst_12.INIT_RAM_1F = 256'h44004240804008168092672208080E0908103020FF4949490001440442444848;
defparam sp_inst_12.INIT_RAM_20 = 256'h242400008047284B00004202A888E98820901010007F15150010000044547F54;
defparam sp_inst_12.INIT_RAM_21 = 256'h92928080FF494949000144044244484890101010020202024202020200222222;
defparam sp_inst_12.INIT_RAM_22 = 256'h9010101080400300030C4080000000E001000000402208044810404080809292;
defparam sp_inst_12.INIT_RAM_23 = 256'h88880000804008168092672208080E0908103020FF4949490001440442444848;
defparam sp_inst_12.INIT_RAM_24 = 256'h101040003F40010E88083010F010FF10080808084126214020106080C80AFF08;
defparam sp_inst_12.INIT_RAM_25 = 256'h92920000402116216710478010F017D8FE02FE0081410D030D11818100101010;
defparam sp_inst_12.INIT_RAM_26 = 256'h44004240001E0202020200002808A8A8A8AC182008080808081E8808E0809292;
defparam sp_inst_12.INIT_RAM_27 = 256'h242400007F89090906010608E628202C22232424007F15150010000044547F54;
defparam sp_inst_12.INIT_RAM_28 = 256'h90004040047F04040404040402F292929292020200FE4242FE00204020222222;
defparam sp_inst_12.INIT_RAM_29 = 256'h56540000000F04040404000000F0101010100000403010102810000016119090;
defparam sp_inst_12.INIT_RAM_2A = 256'h80FEFA02007F000F800000016098808E800780000001460A2222424080005454;
defparam sp_inst_12.INIT_RAM_2B = 256'h04D204D241414040481000000404040400004040475841583F44180820504C50;
defparam sp_inst_12.INIT_RAM_2C = 256'h000000000000000000000000000001010000000000000000000D04D204D204D2;
defparam sp_inst_12.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_13 (
    .DO({sp_inst_13_dout_w[15:0],sp_inst_13_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_13}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_13.READ_MODE = 1'b0;
defparam sp_inst_13.WRITE_MODE = 2'b00;
defparam sp_inst_13.BIT_WIDTH = 16;
defparam sp_inst_13.BLK_SEL = 3'b001;
defparam sp_inst_13.RESET_MODE = "SYNC";
defparam sp_inst_13.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_14 (
    .DO({sp_inst_14_dout_w[15:0],sp_inst_14_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_14}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_14.READ_MODE = 1'b0;
defparam sp_inst_14.WRITE_MODE = 2'b00;
defparam sp_inst_14.BIT_WIDTH = 16;
defparam sp_inst_14.BLK_SEL = 3'b001;
defparam sp_inst_14.RESET_MODE = "SYNC";
defparam sp_inst_14.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_15 (
    .DO({sp_inst_15_dout_w[15:0],sp_inst_15_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_15}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_15.READ_MODE = 1'b0;
defparam sp_inst_15.WRITE_MODE = 2'b00;
defparam sp_inst_15.BIT_WIDTH = 16;
defparam sp_inst_15.BLK_SEL = 3'b001;
defparam sp_inst_15.RESET_MODE = "SYNC";
defparam sp_inst_15.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_16 (
    .DO({sp_inst_16_dout_w[15:0],sp_inst_16_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_16.READ_MODE = 1'b0;
defparam sp_inst_16.WRITE_MODE = 2'b00;
defparam sp_inst_16.BIT_WIDTH = 16;
defparam sp_inst_16.BLK_SEL = 3'b001;
defparam sp_inst_16.RESET_MODE = "SYNC";
defparam sp_inst_16.INIT_RAM_00 = 256'h15005FFF001003AA150003801500028029800010288000100382143850000015;
defparam sp_inst_16.INIT_RAM_01 = 256'h03BF15FF040003BF140004000015040014385FFF028029805800038D15000380;
defparam sp_inst_16.INIT_RAM_02 = 256'h00000000000000004C0006484C00547403BD1500040003800406038814EC0406;
defparam sp_inst_16.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_17 (
    .DO({sp_inst_17_dout_w[15:0],sp_inst_17_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_1}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_17.READ_MODE = 1'b0;
defparam sp_inst_17.WRITE_MODE = 2'b00;
defparam sp_inst_17.BIT_WIDTH = 16;
defparam sp_inst_17.BLK_SEL = 3'b001;
defparam sp_inst_17.RESET_MODE = "SYNC";
defparam sp_inst_17.INIT_RAM_00 = 256'h29BE29BE29BE29BE29BE29BF29BF29BF29BF29BF29BF29BF29BF29BF15000400;
defparam sp_inst_17.INIT_RAM_01 = 256'h440003404400034044000340440003404000036E040029BE29BE29BE29BE29BE;
defparam sp_inst_17.INIT_RAM_02 = 256'h5000549D500054995000549B5000549B5000549B5000549A4400036044000342;
defparam sp_inst_17.INIT_RAM_03 = 256'h28BE28BE28BF28BF28BF28BF28BF28BF28BF28BF28BF15005000549C40000341;
defparam sp_inst_17.INIT_RAM_04 = 256'h2880034004010280298002BF0648040028BE28BE28BE28BE28BE28BE28BE28BE;
defparam sp_inst_17.INIT_RAM_05 = 256'h29BF29BF0280298002BF4C00028028800340040103800280298002BF4C000280;
defparam sp_inst_17.INIT_RAM_06 = 256'h293F001502802980298002BF4C00028028800340298028BF001528BF288028BF;
defparam sp_inst_17.INIT_RAM_07 = 256'h29BE29BE29BE02812981298102BE4C0002802880288003405405157F00152A3F;
defparam sp_inst_17.INIT_RAM_08 = 256'h28BE500029BF29BF28BE500057FF028029BF001128BE640028BE400028BE29BE;
defparam sp_inst_17.INIT_RAM_09 = 256'h28BF29BF002A5C00002128BF28BE293E001002BF28BF0000002A5C00002128BF;
defparam sp_inst_17.INIT_RAM_0A = 256'h600028BF28BF500029BF001500130013001228BF28BF28BE47FF28BF29BF0280;
defparam sp_inst_17.INIT_RAM_0B = 256'h500000670280006728BF6000028028BF29BF00155000283E001002BF02BF28BF;
defparam sp_inst_17.INIT_RAM_0C = 256'h0281288128810015001563FF28BF29BF02BF28BF57FE001500670281006728BF;
defparam sp_inst_17.INIT_RAM_0D = 256'h28BF57FE00152A3F57FE02805C000280283F500029BF02802980298002BF4C00;
defparam sp_inst_17.INIT_RAM_0E = 256'h2980298002BE4C000280288028800015001547FF283F293F2A0028BF29BF0280;
defparam sp_inst_17.INIT_RAM_0F = 256'h500329BF29BF28BF29BF02BF0280298029802980298029802980298029BF0281;
defparam sp_inst_17.INIT_RAM_10 = 256'h02BF2800001028BF028028BF29BF02805C020280283F293F2A00001028BF28BF;
defparam sp_inst_17.INIT_RAM_11 = 256'h28BF29BF028028BF57FE0015288028BF4C002880001002A81C00004068020281;
defparam sp_inst_17.INIT_RAM_12 = 256'h28BF500229BF028028BF29BF028028BF57FD00150067288028BF500229BF0280;
defparam sp_inst_17.INIT_RAM_13 = 256'h0280288028BF500229BF028028BF29BF028028BF57FD001528BF028000152880;
defparam sp_inst_17.INIT_RAM_14 = 256'h28BF02800015288028BF500129BF028028BF29BF028028BF57FC001528BF0280;
defparam sp_inst_17.INIT_RAM_15 = 256'h57FC001528BF02800015288028BF500129BF028028BF29BF028028BF57FC0015;
defparam sp_inst_17.INIT_RAM_16 = 256'h028028BF57FC001528BF02800015288028BF500129BF028028BF29BF028028BF;
defparam sp_inst_17.INIT_RAM_17 = 256'h500029BF29BF028028BF500129BF028028BF57FB0280500129BF028028BF29BF;
defparam sp_inst_17.INIT_RAM_18 = 256'h028028BF29BF028028BF29BF001002BF2800001028BF028028BF001C028028BF;
defparam sp_inst_17.INIT_RAM_19 = 256'h28BF500029BF53FD67FF02802800001028BF028028BF67FD02802800001028BF;
defparam sp_inst_17.INIT_RAM_1A = 256'h28BF028028BF29BF028028BF29BF001002BF2800001028BF028028BF001C0280;
defparam sp_inst_17.INIT_RAM_1B = 256'h5000034057FA028053FD67FF02802800001028BF028028BF67FD028028000010;
defparam sp_inst_17.INIT_RAM_1C = 256'h47FC2800001028BF28BF29BF028028BF57FA00152A3F57FA02805C000280283F;
defparam sp_inst_17.INIT_RAM_1D = 256'h28BF500029BF28BF29BF29BF29BF0280298002BF4C0002812880288000150015;
defparam sp_inst_17.INIT_RAM_1E = 256'h298002BF4C0002802880001528BF47FF29BF02BF28BF2900006728BF29BF0280;
defparam sp_inst_17.INIT_RAM_1F = 256'h02802880034029002A3F28BF43FF034000672A0028BF0340293F001529BF0280;
defparam sp_inst_17.INIT_RAM_20 = 256'h29BF0280298002BF4C0002802880034029800396154A157F0280298002BF4C00;
defparam sp_inst_17.INIT_RAM_21 = 256'h157F00150014001728BF02802881157F440028BF29BF28BF6000028028BF29BF;
defparam sp_inst_17.INIT_RAM_22 = 256'h29BF02BF28BF500029810015157F0015001728BF02802881157F500029810014;
defparam sp_inst_17.INIT_RAM_23 = 256'h02802881157F500029810014157F00150014001728BF02802881157F440028BF;
defparam sp_inst_17.INIT_RAM_24 = 256'h28BF29BF29BF0280298002BF4C0002802880034029810015157F0015001728BF;
defparam sp_inst_17.INIT_RAM_25 = 256'h29810014157F00150014001728BF02802881157F440028BF29BF28BF60000280;
defparam sp_inst_17.INIT_RAM_26 = 256'h440028BF29BF02BF28BF500029810015157F0015001728BF02802881157F5000;
defparam sp_inst_17.INIT_RAM_27 = 256'h001728BF02802881157F500029810014157F00150014001728BF02802881157F;
defparam sp_inst_17.INIT_RAM_28 = 256'h28BF6000028028BF29BF0280298002BF4C0002802880034029810015157F0015;
defparam sp_inst_17.INIT_RAM_29 = 256'h28BF50000015500002805C00001728BF02800014001728BF02802881157F29BF;
defparam sp_inst_17.INIT_RAM_2A = 256'h00150015500002805C00001728BF02800014001728BF02802881157F29BF02BF;
defparam sp_inst_17.INIT_RAM_2B = 256'h4C0002802880034047FF29BF02BF28BF034029BF0280298002BF4C0002802880;
defparam sp_inst_17.INIT_RAM_2C = 256'h288003402900028028BF2900028028BF2980039A140028BF29BF0280298002BF;
defparam sp_inst_17.INIT_RAM_2D = 256'h28BF29BF028029000280157F29BF03A0140329BF29BF0280298002BF4C000280;
defparam sp_inst_17.INIT_RAM_2E = 256'h28BF290002BE157F29000067157F004428BF2900006728BF157F29BF02BF0044;
defparam sp_inst_17.INIT_RAM_2F = 256'h157F400028BF29BF0280298002BF4C0002802880034029000280157F40002A00;
defparam sp_inst_17.INIT_RAM_30 = 256'h400028BF29BF0280298002BF4C0002802880034029000281157F5000290002BE;
defparam sp_inst_17.INIT_RAM_31 = 256'h001502802980298002BF4C00028028800340290002BE157F500029000281157F;
defparam sp_inst_17.INIT_RAM_32 = 256'h0280298002BF4C00028028802880034029000280157F29002A3F157F5400293F;
defparam sp_inst_17.INIT_RAM_33 = 256'h02BF4C0002802880034047FF03402A3F293F2A00157F500029BF293F2A00157F;
defparam sp_inst_17.INIT_RAM_34 = 256'h02BF4C0002802880034029000280157F400003402A3F293F2A00157F02802980;
defparam sp_inst_17.INIT_RAM_35 = 256'h157F298003BA14000380157F2980039014000380157F29800380157F02802980;
defparam sp_inst_17.INIT_RAM_36 = 256'h00200280001C03B228BF29BF0280298002BF4C00028028800340298002800380;
defparam sp_inst_17.INIT_RAM_37 = 256'h00150280298002BF4C0002802880034029800380157F001003BA1400002A5C00;
defparam sp_inst_17.INIT_RAM_38 = 256'h028028800340290000670340157F006700442A3F2900006703402A3F157F293F;
defparam sp_inst_17.INIT_RAM_39 = 256'h00670381157F00672A00157F57FF00152A3F293F001502802980298002BF4C00;
defparam sp_inst_17.INIT_RAM_3A = 256'h28802880034043FF034000672A00157F034043FF034000672A00157F03402900;
defparam sp_inst_17.INIT_RAM_3B = 256'h157F00672A00157F290000670380157F00672A00157F0280298002BF4C000280;
defparam sp_inst_17.INIT_RAM_3C = 256'h0380157F00672A00157F0280298002BF4C0002802880034029000067001402BF;
defparam sp_inst_17.INIT_RAM_3D = 256'h2980298002BF4C00028028800340290000670380157F00672A00157F29000067;
defparam sp_inst_17.INIT_RAM_3E = 256'h02802880288003405454028E1CC700152A3F2900028028821CC7293F00150280;
defparam sp_inst_17.INIT_RAM_3F = 256'h28BF29BF28BF500028BF4400280028BF29BF28BF29BF29BF0280298002BF4C00;

SP sp_inst_18 (
    .DO({sp_inst_18_dout_w[15:0],sp_inst_18_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_2}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_18.READ_MODE = 1'b0;
defparam sp_inst_18.WRITE_MODE = 2'b00;
defparam sp_inst_18.BIT_WIDTH = 16;
defparam sp_inst_18.BLK_SEL = 3'b001;
defparam sp_inst_18.RESET_MODE = "SYNC";
defparam sp_inst_18.INIT_RAM_00 = 256'h280028BF4000280028BF4000280028BF29BF028028BF29BF028028BF500029BF;
defparam sp_inst_18.INIT_RAM_01 = 256'h0015001547FF280028BF29BF028028BF500028BF4400280028BF5BFF280028BF;
defparam sp_inst_18.INIT_RAM_02 = 256'h2A3F157F43FF034000672A00157F0340293F00150280298002BF4C0002802880;
defparam sp_inst_18.INIT_RAM_03 = 256'h57FF028357F628BC1CC70015028602802980298002BF4C000280288003402900;
defparam sp_inst_18.INIT_RAM_04 = 256'h00670044288002BB1CC702802980298002BF4C00028028802880034057FF0280;
defparam sp_inst_18.INIT_RAM_05 = 256'h57FF001500670044288002BA1CC757FF001500670044288002BB1CC757FF0015;
defparam sp_inst_18.INIT_RAM_06 = 256'h001502802980298002BF4C00028028802880034057FE00150067288002BA1CC7;
defparam sp_inst_18.INIT_RAM_07 = 256'h004828BF29BF02802980298002BF4C00028028802880034057FE00152A3F293F;
defparam sp_inst_18.INIT_RAM_08 = 256'h02802980298002BF4C00028028802880034057FE0015006728BF57FE00150067;
defparam sp_inst_18.INIT_RAM_09 = 256'h297F001502802980298002BF4C00028028802880034057FE00152A3F293F0015;
defparam sp_inst_18.INIT_RAM_0A = 256'h02BF4C00028028802880034057FD001500672A7F57FD00150067006F00442A7F;
defparam sp_inst_18.INIT_RAM_0B = 256'h02B41CC7500029BF57FE57FD2900028028B41CC729BF039C1400028029802980;
defparam sp_inst_18.INIT_RAM_0C = 256'h034000672A00157F034067FF028028BF29BF028028BF57FD00152A00001028BF;
defparam sp_inst_18.INIT_RAM_0D = 256'h29000067001502BE157F00672A00157F440028BF29BF02BF28BF500029BF43FF;
defparam sp_inst_18.INIT_RAM_0E = 256'h2A00157F50002900001028BF28B11CC7440028BF43FF034000672A00157F5000;
defparam sp_inst_18.INIT_RAM_0F = 256'h1CC76FFF028028BF29BF028028BF29BF039414002900001028BF28B11CC70067;
defparam sp_inst_18.INIT_RAM_10 = 256'h028002802980298002BF4C00028028802880001502805000001544002A0028B0;
defparam sp_inst_18.INIT_RAM_11 = 256'h29BF2A7F297F001502812980298002BF4C000280288028800015001557FE5413;
defparam sp_inst_18.INIT_RAM_12 = 256'h293F00670044288002AD1CC7293F00670044288002AE1CC7293F0280293F02BF;
defparam sp_inst_18.INIT_RAM_13 = 256'h157F0340293F293F0280293F0067288002AD1CC7293F00670044288002AD1CC7;
defparam sp_inst_18.INIT_RAM_14 = 256'h02BE157F00672A00157F440028BF29BF02BF28BF500029BF43FF034000672A00;
defparam sp_inst_18.INIT_RAM_15 = 256'h2900001028BF28AA1CC7440028BF43FF034000672A00157F5000290000670015;
defparam sp_inst_18.INIT_RAM_16 = 256'h541200152A00001028BF28A91CC72900001028BF28A91CC700672A00157F5000;
defparam sp_inst_18.INIT_RAM_17 = 256'h400028BF29BF57F928A81CC7001502BF6FFF028028BF29BF028028BF29BF2A7F;
defparam sp_inst_18.INIT_RAM_18 = 256'h57FB028057FA57FA02802980298002BF4C0002812880288000150015500028BF;
defparam sp_inst_18.INIT_RAM_19 = 256'h28BF400028BF29BF57FD039C140057FC00152A7F297F028057FB028057FB0280;
defparam sp_inst_18.INIT_RAM_1A = 256'h001502802980298002BF4C0002802880288000152A3F293F02BF5000293F2A00;
defparam sp_inst_18.INIT_RAM_1B = 256'h297F0280006F2A3F57F900152A3F57FB028057FB028057FA028057FA57FA293F;
defparam sp_inst_18.INIT_RAM_1C = 256'h2A3F293F02BF5000293F2A0028BF400028BF29BF57FD039C140057FB00152A7F;
defparam sp_inst_18.INIT_RAM_1D = 256'h028057FA028057FA028057F957F902802980298002BF4C000280288028800015;
defparam sp_inst_18.INIT_RAM_1E = 256'h5000293F2A0028BF400028BF29BF57FC039C140057FA00152A7F297F028057FA;
defparam sp_inst_18.INIT_RAM_1F = 256'h57F9028057F957F802802980298002BF4C0002802880288000152A3F293F02BF;
defparam sp_inst_18.INIT_RAM_20 = 256'h28BF400028BF29BF57FC039C140057FA00152A7F297F028057FA028057F90280;
defparam sp_inst_18.INIT_RAM_21 = 256'h001502802980298002BF4C0002802880288000152A3F293F02BF5000293F2A00;
defparam sp_inst_18.INIT_RAM_22 = 256'h2A7F57F700152A3F57F9028057F9028057F9028057F857F8297F0015293F0015;
defparam sp_inst_18.INIT_RAM_23 = 256'h006F0067006F00442A7F006F2A3F57F7001500672A7F57F700150067006F0044;
defparam sp_inst_18.INIT_RAM_24 = 256'h29BF57FB039C140057F900152A7F297F0280006F0010006F00672A7F006F0010;
defparam sp_inst_18.INIT_RAM_25 = 256'h298002BF4C0002802880288000152A3F293F02BF5000293F2A0028BF400028BF;
defparam sp_inst_18.INIT_RAM_26 = 256'h140057F800152A7F297F028057F8028057F8028057F8028057F757F702802980;
defparam sp_inst_18.INIT_RAM_27 = 256'h02802880288000152A3F293F02BF5000293F2A0028BF400028BF29BF57FA039C;
defparam sp_inst_18.INIT_RAM_28 = 256'h57F657F6297F0015297F0015293F29BF00150015001502802980298002BF4C00;
defparam sp_inst_18.INIT_RAM_29 = 256'h2A7F57F600150067006F00442A7F57F600152A3F57F7028057F7028057F70280;
defparam sp_inst_18.INIT_RAM_2A = 256'h2A7F006F2A3F57F5001500672A7F57F500150067006F00442A7F57F600150067;
defparam sp_inst_18.INIT_RAM_2B = 256'h00672A7F006F0010006F00442A7F006F0010006F00672A7F006F0010006F0044;
defparam sp_inst_18.INIT_RAM_2C = 256'h2A0028BF400028BF29BF57F9039C140057F700152A7F297F0280006F0010006F;
defparam sp_inst_18.INIT_RAM_2D = 256'h28BF294028BF006F0010006F2A00028028BF006F0040006F2A00028028BF293F;
defparam sp_inst_18.INIT_RAM_2E = 256'h293F02BF5000294028BF006F0010006F2A00028028BF006F0040006F2A000280;
defparam sp_inst_18.INIT_RAM_2F = 256'h028002800280542C293F001502802980298002BF4C0002802880288000152A3F;
defparam sp_inst_18.INIT_RAM_30 = 256'h03400340034003400340500029BF03BE1400542F0280028002810280542F0280;
defparam sp_inst_18.INIT_RAM_31 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_18.INIT_RAM_32 = 256'h542B47FF29BF02BF28BF03400340034003400340034003400340034003400340;
defparam sp_inst_18.INIT_RAM_33 = 256'h4C000280288028800340542E0280028002800280542B542F0280028002810280;
defparam sp_inst_18.INIT_RAM_34 = 256'h2A3F4C002880001002911C000040680502802A3F293F293F02802980298002BF;
defparam sp_inst_18.INIT_RAM_35 = 256'h001557F9028044002A3F293F001557F8542E0280028002800280542B293F0280;
defparam sp_inst_18.INIT_RAM_36 = 256'h0280293F542E0281028002810280542E0280028002800280542B44002A3F293F;
defparam sp_inst_18.INIT_RAM_37 = 256'h02800280542A293F02802A3F500457FD00152A3F500457FE00152A3F5004293F;
defparam sp_inst_18.INIT_RAM_38 = 256'h001557F8028044002A3F293F001557F8542D0281028002810280542D02800280;
defparam sp_inst_18.INIT_RAM_39 = 256'h0280293F542D0281028002810280542D0280028002800280542A44002A3F293F;
defparam sp_inst_18.INIT_RAM_3A = 256'h542D02800280028002805429500357FD00152A3F500357FD00152A3F5003293F;
defparam sp_inst_18.INIT_RAM_3B = 256'h542C0280028002800280542944002A3F293F001557F8542D0281028002810280;
defparam sp_inst_18.INIT_RAM_3C = 256'h542C0280028002810280542C02800280028002805429542C0281028002810280;
defparam sp_inst_18.INIT_RAM_3D = 256'h00152A3F542C0280028002810280542C028002800280028054295002293F0280;
defparam sp_inst_18.INIT_RAM_3E = 256'h03400340034003400340034003400340500029BF03BF14005002293F293F57FC;
defparam sp_inst_18.INIT_RAM_3F = 256'h0340034003400340034003400340034003400340034003400340034003400340;

SP sp_inst_19 (
    .DO({sp_inst_19_dout_w[15:0],sp_inst_19_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_3}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_19.READ_MODE = 1'b0;
defparam sp_inst_19.WRITE_MODE = 2'b00;
defparam sp_inst_19.BIT_WIDTH = 16;
defparam sp_inst_19.BLK_SEL = 3'b001;
defparam sp_inst_19.RESET_MODE = "SYNC";
defparam sp_inst_19.INIT_RAM_00 = 256'h2A3F293F001557F747FF29BF02BF28BF03400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_01 = 256'h2A3F293F001554085000293F0280500157FB00152A3F293F5001293F02804400;
defparam sp_inst_19.INIT_RAM_02 = 256'h2A3F680002832A3F293F5C0002802A3F293F02BF2A3F40002A3F293F5C000280;
defparam sp_inst_19.INIT_RAM_03 = 256'h2A3F542E028002800015028002802A3F54270280028002821C000280293F0280;
defparam sp_inst_19.INIT_RAM_04 = 256'h028002800280542744002A3F293F001557F702800015006F2A3F293F5FFF0280;
defparam sp_inst_19.INIT_RAM_05 = 256'h1400542D028002800015028002802A3F54270280028002801C000280542A0280;
defparam sp_inst_19.INIT_RAM_06 = 256'h0340034003400340034003400340034003400340034003400340500029BF03BF;
defparam sp_inst_19.INIT_RAM_07 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_08 = 256'h29BF03BF1400034057F900152A3F293F500047FF29BF02BF28BF034003400340;
defparam sp_inst_19.INIT_RAM_09 = 256'h0340034003400340034003400340034003400340034003400340034003405000;
defparam sp_inst_19.INIT_RAM_0A = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_0B = 256'h298002BF4C00028028802880034053FA580002802A3F47FF29BF02BF28BF0340;
defparam sp_inst_19.INIT_RAM_0C = 256'h001557F3028047FF2A3F293F001557F354280280028002800280542502802980;
defparam sp_inst_19.INIT_RAM_0D = 256'h54500280542544012A3F293F001557F6028000150281001502BF44022A3F293F;
defparam sp_inst_19.INIT_RAM_0E = 256'h0340034003400340034003400340034003400340500029BF03BE1400541F5403;
defparam sp_inst_19.INIT_RAM_0F = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_10 = 256'h03BE1400544F02805403541F47FF29BF02BF28BF034003400340034003400340;
defparam sp_inst_19.INIT_RAM_11 = 256'h03400340034003400340034003400340034003400340034003400340500029BF;
defparam sp_inst_19.INIT_RAM_12 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_13 = 256'h0340500029BF03BF1400541C544F02805423500047FF29BF02BF28BF03400340;
defparam sp_inst_19.INIT_RAM_14 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_15 = 256'h28BF034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_16 = 256'h02BF4C00028028802880034053FD54260280028002800280542347FF29BF02BF;
defparam sp_inst_19.INIT_RAM_17 = 256'h29BF03BF140057F500152A3F5000541B44002A3F293F001557F3028029802980;
defparam sp_inst_19.INIT_RAM_18 = 256'h0340034003400340034003400340034003400340034003400340034003405000;
defparam sp_inst_19.INIT_RAM_19 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_1A = 256'h28BF29BF02802980298002BF4C00028028802880034047FF29BF02BF28BF0340;
defparam sp_inst_19.INIT_RAM_1B = 256'h028028802880034057FF001502802980298002BF4C00028028802880034057E6;
defparam sp_inst_19.INIT_RAM_1C = 256'h02802980298002BF4C00028028802880034057FF028202802980298002BF4C00;
defparam sp_inst_19.INIT_RAM_1D = 256'h002128BF288002A31CC729BF0280298002BF4C00028028802880034057FF0015;
defparam sp_inst_19.INIT_RAM_1E = 256'h2900006728BF157F29000067157F004428BF290002BE157F29BF02BF002A5C00;
defparam sp_inst_19.INIT_RAM_1F = 256'h0340293F00150280298002BF4C0002802880034029000280157F290002BF157F;
defparam sp_inst_19.INIT_RAM_20 = 256'h00150280298002BF4C0002802880034029002A3F157F43FF034000672A00157F;
defparam sp_inst_19.INIT_RAM_21 = 256'h00672A00157F290000670340157F00672A00157F293F02806C0002802A3F293F;
defparam sp_inst_19.INIT_RAM_22 = 256'h2980298002BF4C0002802880034029000067157F00000015000000402A3F0000;
defparam sp_inst_19.INIT_RAM_23 = 256'h28802880034057E00280028057E00280028057E00280028057E0028002800280;
defparam sp_inst_19.INIT_RAM_24 = 256'h03400340034003400340500029BF03A3140057FF02822982298202BD4C000280;
defparam sp_inst_19.INIT_RAM_25 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_26 = 256'h001547FF29BF02BF28BF03400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_27 = 256'h034003400340034003400340500029BF03A314004401001557E0028057DF0280;
defparam sp_inst_19.INIT_RAM_28 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_29 = 256'h0280034047FF29BF02BF28BF0340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_2A = 256'h034003400340034003400340034003400340500029BF03A3140043FF001557DF;
defparam sp_inst_19.INIT_RAM_2B = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_2C = 256'h001557DE02805015028047FF29BF02BF28BF0340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_2D = 256'h03400340034003400340034003400340034003400340500029BF03A314004401;
defparam sp_inst_19.INIT_RAM_2E = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_2F = 256'h03A3140043FF001557DE0280034047FF29BF02BF28BF03400340034003400340;
defparam sp_inst_19.INIT_RAM_30 = 256'h03400340034003400340034003400340034003400340034003400340500029BF;
defparam sp_inst_19.INIT_RAM_31 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_32 = 256'h500029BF03A314004401001557DD02805014028047FF29BF02BF28BF03400340;
defparam sp_inst_19.INIT_RAM_33 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_34 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_35 = 256'h034003400340500029BF03A3140043FF001557DC0280034047FF29BF02BF28BF;
defparam sp_inst_19.INIT_RAM_36 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_37 = 256'h29BF02BF28BF0340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_38 = 256'h03400340034003400340500029BF03A314004401001557DC02805012028047FF;
defparam sp_inst_19.INIT_RAM_39 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_3A = 256'h034047FF29BF02BF28BF03400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_3B = 256'h03400340034003400340034003400340500029BF03A3140043FF001557DB0280;
defparam sp_inst_19.INIT_RAM_3C = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_3D = 256'h001557F95011028047FF29BF02BF28BF03400340034003400340034003400340;
defparam sp_inst_19.INIT_RAM_3E = 256'h034003400340034003400340500029BF03A314004401001557DA028057D90280;
defparam sp_inst_19.INIT_RAM_3F = 256'h0340034003400340034003400340034003400340034003400340034003400340;

SP sp_inst_20 (
    .DO({sp_inst_20_dout_w[15:0],sp_inst_20_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_4}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_20.READ_MODE = 1'b0;
defparam sp_inst_20.WRITE_MODE = 2'b00;
defparam sp_inst_20.BIT_WIDTH = 16;
defparam sp_inst_20.BLK_SEL = 3'b001;
defparam sp_inst_20.RESET_MODE = "SYNC";
defparam sp_inst_20.INIT_RAM_00 = 256'h0280034047FF29BF02BF28BF0340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_01 = 256'h034003400340034003400340034003400340500029BF03A3140043FF001557D9;
defparam sp_inst_20.INIT_RAM_02 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_03 = 256'h001557D90280500F028047FF29BF02BF28BF0340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_04 = 256'h03400340034003400340034003400340034003400340500029BF03A314004401;
defparam sp_inst_20.INIT_RAM_05 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_06 = 256'h03A3140043FF001557D80280034047FF29BF02BF28BF03400340034003400340;
defparam sp_inst_20.INIT_RAM_07 = 256'h03400340034003400340034003400340034003400340034003400340500029BE;
defparam sp_inst_20.INIT_RAM_08 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_09 = 256'h500029BE03A314004401001557D70280500E028047FF29BE02BF28BE03400340;
defparam sp_inst_20.INIT_RAM_0A = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_0B = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_0C = 256'h034003400340500029BE03A3140043FF001557D70280034047FF29BE02BF28BE;
defparam sp_inst_20.INIT_RAM_0D = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_0E = 256'h29BE02BF28BE0340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_0F = 256'h03400340034003400340500029BE03A314004401001557D60280500C028047FF;
defparam sp_inst_20.INIT_RAM_10 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_11 = 256'h034047FF29BE02BF28BE03400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_12 = 256'h03400340034003400340034003400340500029BE03A3140043FF001557D50280;
defparam sp_inst_20.INIT_RAM_13 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_14 = 256'h001557F3500B028047FF29BE02BF28BE03400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_15 = 256'h034003400340034003400340500029BE03A314004401001557D4028057D30280;
defparam sp_inst_20.INIT_RAM_16 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_17 = 256'h0280034047FF29BE02BF28BE0340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_18 = 256'h034003400340034003400340034003400340500029BE03A3140043FF001557D4;
defparam sp_inst_20.INIT_RAM_19 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_1A = 256'h001557D30280500A028047FF29BE02BF28BE0340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_1B = 256'h03400340034003400340034003400340034003400340500029BE03A314004401;
defparam sp_inst_20.INIT_RAM_1C = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_1D = 256'h03A3140043FF001557D20280034047FF29BE02BF28BE03400340034003400340;
defparam sp_inst_20.INIT_RAM_1E = 256'h03400340034003400340034003400340034003400340034003400340500029BE;
defparam sp_inst_20.INIT_RAM_1F = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_20 = 256'h500029BE03A314004401001557D102805008028047FF29BE02BF28BE03400340;
defparam sp_inst_20.INIT_RAM_21 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_22 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_23 = 256'h034003400340500029BE03A3140043FF001557D10280034047FF29BE02BF28BE;
defparam sp_inst_20.INIT_RAM_24 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_25 = 256'h29BE02BF28BE0340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_26 = 256'h03400340034003400340500029BE03A314004401001557D002805007028047FF;
defparam sp_inst_20.INIT_RAM_27 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_28 = 256'h034047FF29BE02BF28BE03400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_29 = 256'h03400340034003400340034003400340500029BE03A3140043FF001557CF0280;
defparam sp_inst_20.INIT_RAM_2A = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_2B = 256'h001557ED5005028047FF29BE02BF28BE03400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_2C = 256'h034003400340034003400340500029BE03A314004401001557CF028057CE0280;
defparam sp_inst_20.INIT_RAM_2D = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_2E = 256'h0280034047FF29BE02BF28BE0340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_2F = 256'h034003400340034003400340034003400340500029BE03A3140043FF001557CE;
defparam sp_inst_20.INIT_RAM_30 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_31 = 256'h001557CD02805004028047FF29BE02BF28BE0340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_32 = 256'h03400340034003400340034003400340034003400340500029BE03A314004401;
defparam sp_inst_20.INIT_RAM_33 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_34 = 256'h03A3140043FF001557CC0280034047FF29BE02BF28BE03400340034003400340;
defparam sp_inst_20.INIT_RAM_35 = 256'h03400340034003400340034003400340034003400340034003400340500029BD;
defparam sp_inst_20.INIT_RAM_36 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_37 = 256'h500029BD03A314004401001557CC02805002028047FF29BD02BF28BD03400340;
defparam sp_inst_20.INIT_RAM_38 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_39 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_3A = 256'h034003400340500029BD03A3140043FF001557CB0280034047FF29BD02BF28BD;
defparam sp_inst_20.INIT_RAM_3B = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_3C = 256'h29BD02BF28BD0340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_3D = 256'h03400340034003400340500029BD03A314004401001557CA02805001028047FF;
defparam sp_inst_20.INIT_RAM_3E = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_20.INIT_RAM_3F = 256'h034047FF29BD02BF28BD03400340034003400340034003400340034003400340;

SP sp_inst_21 (
    .DO({sp_inst_21_dout_w[15:0],sp_inst_21_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_5}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_21.READ_MODE = 1'b0;
defparam sp_inst_21.WRITE_MODE = 2'b00;
defparam sp_inst_21.BIT_WIDTH = 16;
defparam sp_inst_21.BLK_SEL = 3'b001;
defparam sp_inst_21.RESET_MODE = "SYNC";
defparam sp_inst_21.INIT_RAM_00 = 256'h03400340034003400340034003400340500029BD03A3140043FF001557CA0280;
defparam sp_inst_21.INIT_RAM_01 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_21.INIT_RAM_02 = 256'h001500155000028047FF29BD02BF28BD03400340034003400340034003400340;
defparam sp_inst_21.INIT_RAM_03 = 256'h4C00028028802880034057C80280001502802980298002BF4C00028228822882;
defparam sp_inst_21.INIT_RAM_04 = 256'h02802980298002BF4C00028028802880034057C80280028002802980298002BF;
defparam sp_inst_21.INIT_RAM_05 = 256'h034003400340034003400340034003400340500029BF0399140057C702800280;
defparam sp_inst_21.INIT_RAM_06 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_21.INIT_RAM_07 = 256'h0399140057C70280001547FF29BF02BF28BF0340034003400340034003400340;
defparam sp_inst_21.INIT_RAM_08 = 256'h03400340034003400340034003400340034003400340034003400340500029BF;
defparam sp_inst_21.INIT_RAM_09 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_21.INIT_RAM_0A = 256'h034003400340500029BF0399140057C60280028047FF29BF02BF28BF03400340;
defparam sp_inst_21.INIT_RAM_0B = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_21.INIT_RAM_0C = 256'h29BF02BF28BF0340034003400340034003400340034003400340034003400340;
defparam sp_inst_21.INIT_RAM_0D = 256'h57C50280028002802980298002BF4C00028028802880034057C50280001547FF;
defparam sp_inst_21.INIT_RAM_0E = 256'h034003400340034003400340034003400340034003400340500029BF03991400;
defparam sp_inst_21.INIT_RAM_0F = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_21.INIT_RAM_10 = 256'h4C00028028802880034057C50280001547FF29BF02BF28BF0340034003400340;
defparam sp_inst_21.INIT_RAM_11 = 256'h001528BF29BF500029BF02804000001428BF2880157F29BF29BF0280298002BF;
defparam sp_inst_21.INIT_RAM_12 = 256'h2A000380157F2980001528BF157F2880157F29BF0280298002BF4C0002802880;
defparam sp_inst_21.INIT_RAM_13 = 256'h293F001502802980298002BF4C000280288003402900006703800380157F0067;
defparam sp_inst_21.INIT_RAM_14 = 256'h57C5028057C6028057C757C700152A3F57C757C7001557C757C7028157C60280;
defparam sp_inst_21.INIT_RAM_15 = 256'h57C757C6028157C60280293F001502802980298002BF4C000280288028800340;
defparam sp_inst_21.INIT_RAM_16 = 256'h4C00028028802880034057C5028057C6028057C757C600152A3F57C757C60281;
defparam sp_inst_21.INIT_RAM_17 = 256'h03400340034003400340034003400340500029BF0399140002802980298002BF;
defparam sp_inst_21.INIT_RAM_18 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_21.INIT_RAM_19 = 256'h57FE028057FE028247FF29BF02BF28BF03400340034003400340034003400340;
defparam sp_inst_21.INIT_RAM_1A = 256'h57FE028357FE028257FE028157FE028057FE001557FE028357FE028257FE0280;
defparam sp_inst_21.INIT_RAM_1B = 256'h57FD028357FD001557FD028357FE028257FE028057FE028257FE028257FE0282;
defparam sp_inst_21.INIT_RAM_1C = 256'h57FD028257FD028057FD028357FD028057FD028357FD028057FD028357FD0283;
defparam sp_inst_21.INIT_RAM_1D = 256'h28BF29BF29BF02802980298002BF4C00028028802880034057FD028257FD0280;
defparam sp_inst_21.INIT_RAM_1E = 256'h006728BF57FD001500670380006703400067004428BF57FD0015006702BE0067;
defparam sp_inst_21.INIT_RAM_1F = 256'h001502802980298002BF4C00028028802880034057FD00150067038000670340;
defparam sp_inst_21.INIT_RAM_20 = 256'h2A3F500029BF57FC028057FC001557FC0015006702BE006728BF500029BF293F;
defparam sp_inst_21.INIT_RAM_21 = 256'h288003406FFF028028BF29BF028028BF6FFF028128BF29BF028028BF57FD0015;
defparam sp_inst_21.INIT_RAM_22 = 256'h298002BF4C00028028802880034057FF001502802980298002BF4C0002802880;
defparam sp_inst_21.INIT_RAM_23 = 256'h500158010280580002802A3F29BF29BF29BF293F001529BF29BF29BF02802980;
defparam sp_inst_21.INIT_RAM_24 = 256'h57FE28BF28BF29BF028028BF29BF6C00028128BF29BF02BF2A00001028BF28BF;
defparam sp_inst_21.INIT_RAM_25 = 256'h29BF028028BF57FB00152A00001028BF0010001C028028BF02A01C00500029BF;
defparam sp_inst_21.INIT_RAM_26 = 256'h28BF500147FF2A00001028BF28BF29BF028028BF29BF028028BF6FFF028028BF;
defparam sp_inst_21.INIT_RAM_27 = 256'h29BF57FD28BF28BF29BF028028BF29BF6C00028128BF29BF02BF2A00001028BF;
defparam sp_inst_21.INIT_RAM_28 = 256'h028028BF29BF028028BF57FB00152A00001002A61C00001028BF004028BF5000;
defparam sp_inst_21.INIT_RAM_29 = 256'h001002A41C000280001028BF004028BF500029BF57FD28BF0015028028BF6FFF;
defparam sp_inst_21.INIT_RAM_2A = 256'h28BF29BF028028BF29BF028028BF6FFF028028BF29BF028028BF57FA00152A00;
defparam sp_inst_21.INIT_RAM_2B = 256'h29BF29BF02802980298002BF4C000280288028800340034047FE2A00001028BF;
defparam sp_inst_21.INIT_RAM_2C = 256'h2A00001028BF02941CC75000293F57FC28BF28BF29BF00402A3F293F293F0015;
defparam sp_inst_21.INIT_RAM_2D = 256'h57FB28BF0015028028BF6FFF02802A3F293F02802A3F29BF028028BF57FA0015;
defparam sp_inst_21.INIT_RAM_2E = 256'h2A3F293F02802A3F29BF028028BF57F900152A00001028BF02921CC75000293F;
defparam sp_inst_21.INIT_RAM_2F = 256'h29BF29BF29BF29BF29BF02802980298002BF4C0002802880288003406FFF0280;
defparam sp_inst_21.INIT_RAM_30 = 256'h28BF57FE001528BF001500670010006728BF006728BF001028BF004028BF5000;
defparam sp_inst_21.INIT_RAM_31 = 256'h29BF29BF02812980298002BF4C0002802880288003406BFF28BF28BF29BF0280;
defparam sp_inst_21.INIT_RAM_32 = 256'h28BF29BF0280004428BF500029BF004428BF4400034028BF29BF29BF29BF29BF;
defparam sp_inst_21.INIT_RAM_33 = 256'h57F800152A00001028BF29BF028028BF500029BF28BF57FA28BF28BF500029BF;
defparam sp_inst_21.INIT_RAM_34 = 256'h02812880288003406BFF28BF28BF29BF028028BF6BFF28BF28BF29BF028028BF;
defparam sp_inst_21.INIT_RAM_35 = 256'h02BF2A3F29BF29BF293F0015293F0015001529BF29BF02802980298002BF4C00;
defparam sp_inst_21.INIT_RAM_36 = 256'h500029BF57F928BF28BF5C0002802A3F29BF028028BF29BF6C00028128BF29BF;
defparam sp_inst_21.INIT_RAM_37 = 256'h6FFF028028BF29BF028028BF57F700152A00001002971C00001028BF004028BF;
defparam sp_inst_21.INIT_RAM_38 = 256'h2A00001002951C000280001028BF004028BF500029BF57F928BF0015028028BF;
defparam sp_inst_21.INIT_RAM_39 = 256'h028C1C00500029BF57F828BF28BF50006FFF028028BF29BF028028BF57F70015;
defparam sp_inst_21.INIT_RAM_3A = 256'h03406FFF028028BF29BF028028BF57F600152A00001028BF0010001C028028BF;
defparam sp_inst_21.INIT_RAM_3B = 256'h29BF001C28BF28BF500029BF028029BF29BF0280298002BF4C00028028802880;
defparam sp_inst_21.INIT_RAM_3C = 256'h29BF29BF29BF02802980298002BF4C0002802880001528BF47FF29BF02BF28BF;
defparam sp_inst_21.INIT_RAM_3D = 256'h001557FF0280001502BF001128BF2A3F500129BF29BF293F0015293F00150015;
defparam sp_inst_21.INIT_RAM_3E = 256'h6C0028BF001502BF2A3F440028BF29BF002A5C0000210280002A5C00002128BF;
defparam sp_inst_21.INIT_RAM_3F = 256'h57FD001528BF028000152A3F001028BF001C28BF0015006700442A3F440028BF;

SP sp_inst_22 (
    .DO({sp_inst_22_dout_w[15:0],sp_inst_22_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_6}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_22.READ_MODE = 1'b0;
defparam sp_inst_22.WRITE_MODE = 2'b00;
defparam sp_inst_22.BIT_WIDTH = 16;
defparam sp_inst_22.BLK_SEL = 3'b001;
defparam sp_inst_22.RESET_MODE = "SYNC";
defparam sp_inst_22.INIT_RAM_00 = 256'h2A3F00670280006728BF001028BF001C28BF0015006700442A3F29BF02805000;
defparam sp_inst_22.INIT_RAM_01 = 256'h4C0002802880288003406BFE28BF2A3F29BF028028BF57FC001528BF00150015;
defparam sp_inst_22.INIT_RAM_02 = 256'h57B70280028057B70280028057B70280028057B70280028002802980298002BF;
defparam sp_inst_22.INIT_RAM_03 = 256'h001557B70280028057B70280028057B70280028057B70280028057B702800280;
defparam sp_inst_22.INIT_RAM_04 = 256'h0280001557B60280001557B70280001557B70280001557B70280028057B70280;
defparam sp_inst_22.INIT_RAM_05 = 256'h03400340034003400340034003400340034003400340500029BF03BF140057B6;
defparam sp_inst_22.INIT_RAM_06 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_07 = 256'h028057B70280028057B70280028047FF29BF02BF28BF03400340034003400340;
defparam sp_inst_22.INIT_RAM_08 = 256'h2880034057B60280001557B70280028057B70280028057B70280028057B70280;
defparam sp_inst_22.INIT_RAM_09 = 256'h29BF0399140057B8001502BF57B8001502BF02802980298002BF4C0002802880;
defparam sp_inst_22.INIT_RAM_0A = 256'h0340034003400340034003400340034003400340034003400340034003405000;
defparam sp_inst_22.INIT_RAM_0B = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_0C = 256'h140057BA02802980298002BF4C00028028802880034047FF29BF02BF28BF0340;
defparam sp_inst_22.INIT_RAM_0D = 256'h0340034003400340034003400340034003400340034003400340500029BF0399;
defparam sp_inst_22.INIT_RAM_0E = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_0F = 256'h02802980298002BF4C00028028802880034047FF29BF02BF28BF034003400340;
defparam sp_inst_22.INIT_RAM_10 = 256'h57BF540057F457F157D202802980298002BF4C00028028802880034057BA0280;
defparam sp_inst_22.INIT_RAM_11 = 256'h034003400340500029BF0399140002802980298002BF4C000280288028800340;
defparam sp_inst_22.INIT_RAM_12 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_13 = 256'h29BF02BF28BF0340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_14 = 256'h0340034003400340034003400340034003400340500029BF03911400540547FF;
defparam sp_inst_22.INIT_RAM_15 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_16 = 256'h0340500029BF03911400540547FF29BF02BF28BF034003400340034003400340;
defparam sp_inst_22.INIT_RAM_17 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_18 = 256'h28BF034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_19 = 256'h03400340034003400340034003400340500029BF03911400540847FF29BF02BF;
defparam sp_inst_22.INIT_RAM_1A = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_1B = 256'h288028800340540647FF29BF02BF28BF03400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_1C = 256'h001502BE00000341000000402A3F293F293F001502802980298002BF4C000280;
defparam sp_inst_22.INIT_RAM_1D = 256'h00672A00157F034043FF034000672A00157F034029002A3F157F57B7293F0000;
defparam sp_inst_22.INIT_RAM_1E = 256'h2A00157F034043FF034000672A00157F03402900157F293F2A00157F47FF0340;
defparam sp_inst_22.INIT_RAM_1F = 256'h034003400340034003400340500029BF028057B7293F2A00157F47FF03400067;
defparam sp_inst_22.INIT_RAM_20 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_21 = 256'h00152A3F47FF29BF02BF28BF0340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_22 = 256'h006700402A3F293F0015293F0015001502802980298002BF4C00028028802880;
defparam sp_inst_22.INIT_RAM_23 = 256'h00672A00157F034043FF034000672A00157F034029002A3F157F57B6293F0341;
defparam sp_inst_22.INIT_RAM_24 = 256'h157F034043FF034000672A00157F034029002A3F157F293F2A00157F47FF0340;
defparam sp_inst_22.INIT_RAM_25 = 256'h03400340034003400340500029BF028057B5293F2A00157F47FF034000672A00;
defparam sp_inst_22.INIT_RAM_26 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_27 = 256'h034047FF29BF02BF28BF03400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_28 = 256'h00152A3F293F293F0015293F0015001502802980298002BF4C00028028802880;
defparam sp_inst_22.INIT_RAM_29 = 256'h028028802880034057FE001500152A3F0067000000152A3F283F293F001557FC;
defparam sp_inst_22.INIT_RAM_2A = 256'h293F001557FC00152A3F293F293F0015293F0015001502802980298002BF4C00;
defparam sp_inst_22.INIT_RAM_2B = 256'h4C00028028802880034057FD001500152A3F0067000000142A3F00000014283F;
defparam sp_inst_22.INIT_RAM_2C = 256'h034003400340034003400340500029BF028B57AE0280028002802980298002BF;
defparam sp_inst_22.INIT_RAM_2D = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_2E = 256'h0280001547FF29BF02BF28BF0340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_2F = 256'h034003400340034003400340034003400340034003400340500029BF028B57AD;
defparam sp_inst_22.INIT_RAM_30 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_31 = 256'h29BF028B57FC0280028057AC0280028047FF29BF02BF28BF0340034003400340;
defparam sp_inst_22.INIT_RAM_32 = 256'h0340034003400340034003400340034003400340034003400340034003405000;
defparam sp_inst_22.INIT_RAM_33 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_34 = 256'h0280028257FB0280001557FB0280028057FB0280028047FF29BF02BF28BF0340;
defparam sp_inst_22.INIT_RAM_35 = 256'h2980298002BF4C000280288028800015001557FB0280028157FB0280028057FB;
defparam sp_inst_22.INIT_RAM_36 = 256'h034003400340034003400340034003400340500029BF028E57FB028002810280;
defparam sp_inst_22.INIT_RAM_37 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_38 = 256'h2A3F293F001557F8028047FF29BF02BF28BF0340034003400340034003400340;
defparam sp_inst_22.INIT_RAM_39 = 256'h298002BF4C000280288028800340293F001557F8028057FB0280028044000340;
defparam sp_inst_22.INIT_RAM_3A = 256'h0015028029802980298002BF4C00028028802880034057FB0280028002802980;
defparam sp_inst_22.INIT_RAM_3B = 256'h5C000280580002802A3F293F293F293F02BF293F0015293F29BF29BF001529BF;
defparam sp_inst_22.INIT_RAM_3C = 256'h00150067001502BE2A3F03405000293F0280293F02815000293F0280293F0280;
defparam sp_inst_22.INIT_RAM_3D = 256'h001028BF28BF500029BF57FA0280028257F90280001557FB0280028257F90280;
defparam sp_inst_22.INIT_RAM_3E = 256'h02802A3F57F8028000152A3F63FF28BF2A3F29BF028028BF57F9028000152A00;
defparam sp_inst_22.INIT_RAM_3F = 256'h400028BF29BF02BF28BF293F001557F7028029BF03A2140057FA028002825C00;

SP sp_inst_23 (
    .DO({sp_inst_23_dout_w[15:0],sp_inst_23_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_7}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_23.READ_MODE = 1'b0;
defparam sp_inst_23.WRITE_MODE = 2'b00;
defparam sp_inst_23.BIT_WIDTH = 16;
defparam sp_inst_23.BLK_SEL = 3'b001;
defparam sp_inst_23.RESET_MODE = "SYNC";
defparam sp_inst_23.INIT_RAM_00 = 256'h001557F60280400128BF57FA0280028243FF006700142A3F2A3F440003402A3F;
defparam sp_inst_23.INIT_RAM_01 = 256'h57F602805C0002802A3F293F02BF40000340006700142A3F2A3F293F44000340;
defparam sp_inst_23.INIT_RAM_02 = 256'h298028BF00102A3F004002BF2A3F40002A3F293F0340001557F60280293F0015;
defparam sp_inst_23.INIT_RAM_03 = 256'h500029BF293F02806C0002802A3F293F028044002A3F298028BF00402A3F5000;
defparam sp_inst_23.INIT_RAM_04 = 256'h293F02BF500063FF28BF2A3F29BF028028BF2900001557F50280001028BF28BF;
defparam sp_inst_23.INIT_RAM_05 = 256'h2980298002BF4C0002802880288028800015283F57F70280001557F802800282;
defparam sp_inst_23.INIT_RAM_06 = 256'h02BF293F2A3F57F80280028057F60280028057F802800280293F29BF00150281;
defparam sp_inst_23.INIT_RAM_07 = 256'h2A3F5C00028028BF4400283F293F001557FC0280001502800015001502BF02BF;
defparam sp_inst_23.INIT_RAM_08 = 256'h02BF4C000281288028800015283F293F02BF500029002A3F028028BF290028BF;
defparam sp_inst_23.INIT_RAM_09 = 256'h293F02BE57F80280028257F60280001557F802800280293F29BF028129802980;
defparam sp_inst_23.INIT_RAM_0A = 256'h293F4400283F293F001557FC0280001502800015001502BF02BF02BF293F0280;
defparam sp_inst_23.INIT_RAM_0B = 256'h293F00152A3F2A3F001002BF2A3F29002A3F001002BF001028BF2A3F2A3F5000;
defparam sp_inst_23.INIT_RAM_0C = 256'h02800282293F02BF58002A3F2A3F001002BF2A3F6FFF02802A3F293F02802A3F;
defparam sp_inst_23.INIT_RAM_0D = 256'h57FD028128B21CC7297F02802980298002BF4C000281288028800015283F57F6;
defparam sp_inst_23.INIT_RAM_0E = 256'h006F001C0280006F006700442A0028B11CC74400001557FE28B21CC744000015;
defparam sp_inst_23.INIT_RAM_0F = 256'h298002BF4C0002802880288000152A7F297F0010006F0340006F2A0028B11CC7;
defparam sp_inst_23.INIT_RAM_10 = 256'h298028BF0280288028BF29002A3F0010288028BF288028BF293F001529BF0280;
defparam sp_inst_23.INIT_RAM_11 = 256'h288028BF288028BF298028BF0280288028BF298028BF6000288028BF288028BF;
defparam sp_inst_23.INIT_RAM_12 = 256'h28BF6000288028BF288028BF298028BF0280288028BF298028BF288028BF6400;
defparam sp_inst_23.INIT_RAM_13 = 256'h57C20384140057EF57ED57EE57EB02802980298002BF4C000280288003402980;
defparam sp_inst_23.INIT_RAM_14 = 256'h034003400340034003400340034003400340034003400340500029BF03BF1400;
defparam sp_inst_23.INIT_RAM_15 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_23.INIT_RAM_16 = 256'h034003400340500029BF03BF140057EE47FF29BF02BF28BF0340034003400340;
defparam sp_inst_23.INIT_RAM_17 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_23.INIT_RAM_18 = 256'h29BF02BF28BF0340034003400340034003400340034003400340034003400340;
defparam sp_inst_23.INIT_RAM_19 = 256'h290002B31CC70015001557C257DA290002B41CC75C0C0280001557A3028047FF;
defparam sp_inst_23.INIT_RAM_1A = 256'h5C0002802A00028F1CC74C002880001002911C000040680C02802A0002901CC7;
defparam sp_inst_23.INIT_RAM_1B = 256'h028E1CC729000280028E1CC75C0002802A0002B21CC72900028F1CC7540D0280;
defparam sp_inst_23.INIT_RAM_1C = 256'h29000280028D1CC729000280028D1CC75C0C02802A0002B11CC7500C29000280;
defparam sp_inst_23.INIT_RAM_1D = 256'h5C0002802A0002AF1CC72900028C1CC7540C02805C0002802A00028D1CC7500C;
defparam sp_inst_23.INIT_RAM_1E = 256'h028B1CC75C0002802A0002AF1CC7500B29000280028C1CC729000280028C1CC7;
defparam sp_inst_23.INIT_RAM_1F = 256'h29000280028A1CC75C0002802A0002AE1CC7500B29000280028B1CC729000280;
defparam sp_inst_23.INIT_RAM_20 = 256'h02891CC72900028002891CC75C0B02802A0002AD1CC7500B29000280028A1CC7;
defparam sp_inst_23.INIT_RAM_21 = 256'h02AB1CC75417290002881CC7540B02805C0002802A0002891CC7500B29000280;
defparam sp_inst_23.INIT_RAM_22 = 256'h02802A0002871CC7500A2900028002871CC72900028002881CC75C0A02802A00;
defparam sp_inst_23.INIT_RAM_23 = 256'h2900028002861CC75C0A02802A0002AA1CC75419290002871CC7540B02805C00;
defparam sp_inst_23.INIT_RAM_24 = 256'h1CC7290002851CC7540A02805C0002802A0002861CC7500A2900028002861CC7;
defparam sp_inst_23.INIT_RAM_25 = 256'h2A0002A71CC7500A2900028002841CC72900028002851CC75C0002802A0002A8;
defparam sp_inst_23.INIT_RAM_26 = 256'h5C0002802A0002A61CC750092900028002841CC72900028002841CC75C000280;
defparam sp_inst_23.INIT_RAM_27 = 256'h02821CC75C0902802A0002A61CC750092900028002831CC72900028002831CC7;
defparam sp_inst_23.INIT_RAM_28 = 256'h02811CC7540902805C0002802A0002811CC750092900028002821CC729000280;
defparam sp_inst_23.INIT_RAM_29 = 256'h1CC750092900028002801CC72900028002811CC75C0002802A0002A41CC72900;
defparam sp_inst_23.INIT_RAM_2A = 256'h2A0002A21CC750082900028002BF1CC72900028002801CC75C0002802A0002A3;
defparam sp_inst_23.INIT_RAM_2B = 256'h5C0802802A0002A11CC750082900028002BF1CC72900028002BF1CC75C000280;
defparam sp_inst_23.INIT_RAM_2C = 256'h540802805C0002802A0002BD1CC750082900028002BE1CC72900028002BE1CC7;
defparam sp_inst_23.INIT_RAM_2D = 256'h2900028002BC1CC72900028002BC1CC75C0002802A0002A01CC7290002BD1CC7;
defparam sp_inst_23.INIT_RAM_2E = 256'h1CC750072900028002BB1CC72900028002BC1CC75C0002802A00029F1CC75008;
defparam sp_inst_23.INIT_RAM_2F = 256'h2A00029D1CC750072900028002BA1CC72900028002BB1CC75C0002802A00029E;
defparam sp_inst_23.INIT_RAM_30 = 256'h5C0002802A0002B91CC750072900028002BA1CC72900028002BA1CC75C070280;
defparam sp_inst_23.INIT_RAM_31 = 256'h1CC72900028002B81CC75C0702802A00029C1CC7541B290002B91CC754070280;
defparam sp_inst_23.INIT_RAM_32 = 256'h1CC7540F290002B71CC7540702805C0002802A0002B81CC750072900028002B8;
defparam sp_inst_23.INIT_RAM_33 = 256'h2A0002B61CC750062900028002B61CC72900028002B71CC75C0602802A00029A;
defparam sp_inst_23.INIT_RAM_34 = 256'h028002B51CC75C0602802A0002991CC7541F290002B61CC7540602805C000280;
defparam sp_inst_23.INIT_RAM_35 = 256'h290002B41CC7540602805C0002802A0002B51CC750062900028002B51CC72900;
defparam sp_inst_23.INIT_RAM_36 = 256'h02961CC750052900028002B31CC72900028002B41CC75C0002802A0002971CC7;
defparam sp_inst_23.INIT_RAM_37 = 256'h02802A0002951CC750052900028002B21CC72900028002B31CC75C0002802A00;
defparam sp_inst_23.INIT_RAM_38 = 256'h02805C0002802A0002B11CC750052900028002B21CC72900028002B21CC75C05;
defparam sp_inst_23.INIT_RAM_39 = 256'h02B01CC72900028002B01CC75C0502802A0002941CC7290002B11CC754215405;
defparam sp_inst_23.INIT_RAM_3A = 256'h2A0002921CC7290002AF1CC7540502805C0002802A0002B01CC7500529000280;
defparam sp_inst_23.INIT_RAM_3B = 256'h5C0002802A0002911CC750042900028002AF1CC72900028002AF1CC75C000280;
defparam sp_inst_23.INIT_RAM_3C = 256'h02AD1CC75C0402802A0002911CC750042900028002AE1CC72900028002AE1CC7;
defparam sp_inst_23.INIT_RAM_3D = 256'h1CC7540F540402805C0002802A0002AC1CC750042900028002AD1CC729000280;
defparam sp_inst_23.INIT_RAM_3E = 256'h50042900028002AB1CC72900028002AB1CC75C0402802A00028F1CC7290002AC;
defparam sp_inst_23.INIT_RAM_3F = 256'h57B22900028002AA1CC72900028002AA1CC7540402805C0002802A0002AB1CC7;

SP sp_inst_24 (
    .DO({sp_inst_24_dout_w[15:0],sp_inst_24_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_8}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_24.READ_MODE = 1'b0;
defparam sp_inst_24.WRITE_MODE = 2'b00;
defparam sp_inst_24.BIT_WIDTH = 16;
defparam sp_inst_24.BLK_SEL = 3'b001;
defparam sp_inst_24.RESET_MODE = "SYNC";
defparam sp_inst_24.INIT_RAM_00 = 256'h02A91CC750032900028002A91CC72900028002AA1CC75C0302802A00028D1CC7;
defparam sp_inst_24.INIT_RAM_01 = 256'h028002A81CC75C0002802A00028C1CC7290002A91CC7540302805C0002802A00;
defparam sp_inst_24.INIT_RAM_02 = 256'h1CC72900028002A71CC75C0002802A00028B1CC750032900028002A81CC72900;
defparam sp_inst_24.INIT_RAM_03 = 256'h028002A61CC72900028002A61CC75C0002802A00028A1CC750032900028002A7;
defparam sp_inst_24.INIT_RAM_04 = 256'h50022900028002A51CC72900028002A51CC75C0202802A0002891CC750022900;
defparam sp_inst_24.INIT_RAM_05 = 256'h57AB2900028002A41CC72900028002A41CC7540202805C0002802A0002A51CC7;
defparam sp_inst_24.INIT_RAM_06 = 256'h02A31CC750022900028002A31CC72900028002A41CC75C0202802A0002871CC7;
defparam sp_inst_24.INIT_RAM_07 = 256'h028002A21CC75C0002802A0002861CC7290002A31CC7540202805C0002802A00;
defparam sp_inst_24.INIT_RAM_08 = 256'h1CC72900028002A11CC75C0002802A0002851CC750012900028002A21CC72900;
defparam sp_inst_24.INIT_RAM_09 = 256'h028002A01CC72900028002A01CC75C0102802A0002841CC750012900028002A1;
defparam sp_inst_24.INIT_RAM_0A = 256'h029F1CC729000280029F1CC757B3540102805C0002802A0002A01CC750012900;
defparam sp_inst_24.INIT_RAM_0B = 256'h500029000280029E1CC729000280029E1CC75C0102802A0002821CC729000280;
defparam sp_inst_24.INIT_RAM_0C = 256'h029D1CC729000280029D1CC757CD2900028002811CC757D544002A0002811CC7;
defparam sp_inst_24.INIT_RAM_0D = 256'h034053F2034053F2034053F2034053F2034053F2034053F2034053F229000280;
defparam sp_inst_24.INIT_RAM_0E = 256'h034053F2034053F2034053F2034053F2034053F2034053F2034053F2034053F2;
defparam sp_inst_24.INIT_RAM_0F = 256'h001502802980298002BF53F2034053F2034053F2034053F2034053F2034053F2;
defparam sp_inst_24.INIT_RAM_10 = 256'h00150281028002951C0057D44C0028800010029D1C000040680802802A7F297F;
defparam sp_inst_24.INIT_RAM_11 = 256'h0280028057D602810280028057D602800280028057D600150280028057D80280;
defparam sp_inst_24.INIT_RAM_12 = 256'h028057D402800280029A1C00028057D7028000150280028057D4500857D60281;
defparam sp_inst_24.INIT_RAM_13 = 256'h028057D6028002800280028057D302800280029A1C00028057D7028002800280;
defparam sp_inst_24.INIT_RAM_14 = 256'h500757D6028102800280028057D6028002800280028057D30280028002991C00;
defparam sp_inst_24.INIT_RAM_15 = 256'h0280028002971C00028057D6028100150280028057D6028000150280028057D3;
defparam sp_inst_24.INIT_RAM_16 = 256'h57D20280028002961C00028057D6028002800280028057D502800280028057D3;
defparam sp_inst_24.INIT_RAM_17 = 256'h57D20280028002951C00028057D5028102800280028057D60280028002800280;
defparam sp_inst_24.INIT_RAM_18 = 256'h57D402800015028057D2500657D5028102800280028057D50280028002800280;
defparam sp_inst_24.INIT_RAM_19 = 256'h500657D5001502800280028057D5028000150280028057D50280001502800280;
defparam sp_inst_24.INIT_RAM_1A = 256'h02800281028057D1500557D5001502800280028057D5028000150280028057D2;
defparam sp_inst_24.INIT_RAM_1B = 256'h0280028057D4001500150280028057D1500557D5028102800280028057D50280;
defparam sp_inst_24.INIT_RAM_1C = 256'h028057D1500557D4001502800280028057D4028100150280028057D402800015;
defparam sp_inst_24.INIT_RAM_1D = 256'h0280028057D1500557D302810280028057D302810280028057D4028002800281;
defparam sp_inst_24.INIT_RAM_1E = 256'h1C00028057D4028000150280028057D302800015028057D0500457D402800280;
defparam sp_inst_24.INIT_RAM_1F = 256'h028D1C00028057D202810280028057D3028002800280028057D002800280028E;
defparam sp_inst_24.INIT_RAM_20 = 256'h57D202810280028057D202810280028057D3028002800280028057D002800280;
defparam sp_inst_24.INIT_RAM_21 = 256'h00150280028057D0500457D3028002800280028057D002800280028C1C000280;
defparam sp_inst_24.INIT_RAM_22 = 256'h02800280028057D002800280028A1C00028057D3028100150280028057D30280;
defparam sp_inst_24.INIT_RAM_23 = 256'h02800280028057CF0280028002891C00028057D3028102800280028057D30280;
defparam sp_inst_24.INIT_RAM_24 = 256'h0280028002881C00028057D102810280028057D2028102800280028057D20280;
defparam sp_inst_24.INIT_RAM_25 = 256'h02810015028057D2028000150280028057CF500357D2028002800280028057CF;
defparam sp_inst_24.INIT_RAM_26 = 256'h028057CE500257D2028100150280028057D2028000150280028057CF500357D1;
defparam sp_inst_24.INIT_RAM_27 = 256'h028057D1028002800280028057CE500257D2028002800280028057D102800280;
defparam sp_inst_24.INIT_RAM_28 = 256'h0015028057D1028000150280028057CE500257D002810280028057D002800280;
defparam sp_inst_24.INIT_RAM_29 = 256'h57CE500257D002810280028057D000150280028057D002810015028057D00281;
defparam sp_inst_24.INIT_RAM_2A = 256'h0280028057D002810280028057D1028002800280028057D10280028002800280;
defparam sp_inst_24.INIT_RAM_2B = 256'h02800280028057D0028002800280028057CD500157D002810280028057D00015;
defparam sp_inst_24.INIT_RAM_2C = 256'h1C00028057D0028100150280028057D0028000150280028057CD500157D00280;
defparam sp_inst_24.INIT_RAM_2D = 256'h1C00028057D0028102800280028057D0028002800280028057CD028002800280;
defparam sp_inst_24.INIT_RAM_2E = 256'h0280028057D0028102800280028057D0028002800280028057CD0280028002BF;
defparam sp_inst_24.INIT_RAM_2F = 256'h028057CC500057CF028002800280028057CC0280028002BE1C00028057CF0281;
defparam sp_inst_24.INIT_RAM_30 = 256'h00150280028057CE02810280028057CF028002800280028057CF028002800280;
defparam sp_inst_24.INIT_RAM_31 = 256'h028100150280028057CF028000150280028057CC500057CE02810280028057CE;
defparam sp_inst_24.INIT_RAM_32 = 256'h40012A7F297F001557E602802980298002BF4C000280288028800340034057CF;
defparam sp_inst_24.INIT_RAM_33 = 256'h29800010004028BF02B61CC728800010004002B61CC702BF28BF500029BF0280;
defparam sp_inst_24.INIT_RAM_34 = 256'h57D1028002800015028002802A7F298002B51CC72A7F63FF28BF29BF02BF28BF;
defparam sp_inst_24.INIT_RAM_35 = 256'h034003400340034003400340034003400340034003400340500029BF03BF1400;
defparam sp_inst_24.INIT_RAM_36 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_24.INIT_RAM_37 = 256'h0340500029BF03B2140057C357F6028047FF29BF02BF28BF0340034003400340;
defparam sp_inst_24.INIT_RAM_38 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_24.INIT_RAM_39 = 256'h28BF034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_24.INIT_RAM_3A = 256'h4C0002802880288003402900028002AF1CC72900028002B01CC747FF29BF02BF;
defparam sp_inst_24.INIT_RAM_3B = 256'h28BF29BF028028BF29800010004028BF02AE1CC7500029BF02802980298002BF;
defparam sp_inst_24.INIT_RAM_3C = 256'h034003400340034003400340034003400340500029BF03B2140057C26FFF0280;
defparam sp_inst_24.INIT_RAM_3D = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_24.INIT_RAM_3E = 256'h1CC72900028002AB1CC747FF29BF02BF28BF0340034003400340034003400340;
defparam sp_inst_24.INIT_RAM_3F = 256'h2A7F297F001557E302802980298002BF4C0002802880288003402900028002AB;

SP sp_inst_25 (
    .DO({sp_inst_25_dout_w[15:0],sp_inst_25_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_9}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_25.READ_MODE = 1'b0;
defparam sp_inst_25.WRITE_MODE = 2'b00;
defparam sp_inst_25.BIT_WIDTH = 16;
defparam sp_inst_25.BLK_SEL = 3'b001;
defparam sp_inst_25.RESET_MODE = "SYNC";
defparam sp_inst_25.INIT_RAM_00 = 256'h57A657F302805C0128800010004028BF02A91CC72A7F6802028028BF29BF4002;
defparam sp_inst_25.INIT_RAM_01 = 256'h03400340034003400340034003400340034003400340500029BF03BE140057C3;
defparam sp_inst_25.INIT_RAM_02 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_03 = 256'h29BF03BE140057F2028057A657C247FF29BF02BF28BF03400340034003400340;
defparam sp_inst_25.INIT_RAM_04 = 256'h0340034003400340034003400340034003400340034003400340034003405000;
defparam sp_inst_25.INIT_RAM_05 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_06 = 256'h57F2028050002900028002A31CC72900028002A41CC747FF29BF02BF28BF0340;
defparam sp_inst_25.INIT_RAM_07 = 256'h03400340034003400340034003400340034003400340500029BF03BF140057BF;
defparam sp_inst_25.INIT_RAM_08 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_09 = 256'h0280288028800340034057F1028047FF29BF02BF28BF03400340034003400340;
defparam sp_inst_25.INIT_RAM_0A = 256'h1CC7680202802A0002831CC740052A0002831CC729BF02802980298002BF4C00;
defparam sp_inst_25.INIT_RAM_0B = 256'h02802A0002811CC7298028B41CC7001C0280288028B51CC768000280288028B5;
defparam sp_inst_25.INIT_RAM_0C = 256'h0280288028B31CC7298028B31CC70010288028B41CC700150067002A5C000021;
defparam sp_inst_25.INIT_RAM_0D = 256'h0021028028BF500029BF02BF288028B21CC729BF288028B31CC7298028B31CC7;
defparam sp_inst_25.INIT_RAM_0E = 256'h028028BF028002800280004028BF29BF002A5C000021028028BF29BF002A5C00;
defparam sp_inst_25.INIT_RAM_0F = 256'h03400340034003400340500029BF03B3140067FF28BF29BF02BF28BF57CB0015;
defparam sp_inst_25.INIT_RAM_10 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_11 = 256'h29BF47FF29BF02BF28BF03400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_12 = 256'h028028BF57C400150280029A1C00028002800040001128BF288028AE1CC75000;
defparam sp_inst_25.INIT_RAM_13 = 256'h28AC1CC728800010004028BF02961CC7500029BF6BFF288028AD1CC728BF29BF;
defparam sp_inst_25.INIT_RAM_14 = 256'h5C0202802A0002B81CC76FFF028028BF29BF028028BF500029BF02805C002880;
defparam sp_inst_25.INIT_RAM_15 = 256'h034003400340034003400340500029BF03BE140057BE57A157EE0280400128BF;
defparam sp_inst_25.INIT_RAM_16 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_17 = 256'h57A157BD47FF29BF02BF28BF0340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_18 = 256'h0340034003400340034003400340034003400340500029BF03BE140057ED0280;
defparam sp_inst_25.INIT_RAM_19 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_1A = 256'h028F1CC729000280028F1CC747FF29BF02BF28BF034003400340034003400340;
defparam sp_inst_25.INIT_RAM_1B = 256'h29BF03BF140057A057BA57ED02805000298028A41CC7298028A51CC729000280;
defparam sp_inst_25.INIT_RAM_1C = 256'h0340034003400340034003400340034003400340034003400340034003405000;
defparam sp_inst_25.INIT_RAM_1D = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_1E = 256'h2A0002AE1CC757EC0280298028A11CC7298028A21CC747FF29BF02BF28BF0340;
defparam sp_inst_25.INIT_RAM_1F = 256'h028D1C0002800280004028BF500029BF298028A01CC7298028A11CC75C000280;
defparam sp_inst_25.INIT_RAM_20 = 256'h298002BF4C00028028802880034067FF028028BF29BF028028BF57C000150280;
defparam sp_inst_25.INIT_RAM_21 = 256'h680002802880289E1CC7680102802A0002AC1CC740042A0002AC1CC702802980;
defparam sp_inst_25.INIT_RAM_22 = 256'h0067002A5C00002102802A0002AB1CC72980289E1CC7001C02802880289E1CC7;
defparam sp_inst_25.INIT_RAM_23 = 256'h1CC72980289C1CC702802880289C1CC72980289D1CC700102880289D1CC70015;
defparam sp_inst_25.INIT_RAM_24 = 256'h28BF293F002A5C000020028028BF500029BF02BF2880289B1CC729BF2880289C;
defparam sp_inst_25.INIT_RAM_25 = 256'h57C500150280001502800280283F00150280004028BF29BF002A5C0000200280;
defparam sp_inst_25.INIT_RAM_26 = 256'h0340034003400340034003400340500029BF03A6140067FF28BF29BF02BF28BF;
defparam sp_inst_25.INIT_RAM_27 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_28 = 256'h2A0002A41CC747FF29BF02BF28BF034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_29 = 256'h028002801CC72900028002801CC757E902805C000291288028971CC75C010280;
defparam sp_inst_25.INIT_RAM_2A = 256'h03400340034003400340034003400340034003400340500029BF03BF14002900;
defparam sp_inst_25.INIT_RAM_2B = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_2C = 256'h5000298028931CC7298028931CC747FF29BF02BF28BF03400340034003400340;
defparam sp_inst_25.INIT_RAM_2D = 256'h03400340034003400340034003400340500029BF03BF140057B557E8028057BD;
defparam sp_inst_25.INIT_RAM_2E = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_2F = 256'h2900028002BA1CC747FF29BF02BF28BF03400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_30 = 256'h1CC75C0002802A00029D1CC72980288F1CC7298028901CC72900028002BA1CC7;
defparam sp_inst_25.INIT_RAM_31 = 256'h57BC0015028002BB1C0002800280004028BF500029BF2980288F1CC72980288F;
defparam sp_inst_25.INIT_RAM_32 = 256'h1CC702802980298002BF4C00028028802880034067FF028028BF29BF028028BF;
defparam sp_inst_25.INIT_RAM_33 = 256'h2880288C1CC7680002802880288C1CC7680102802A00029A1CC740032A00029A;
defparam sp_inst_25.INIT_RAM_34 = 256'h288B1CC700150067002A5C00002102802A0002991CC72980288C1CC7001C0280;
defparam sp_inst_25.INIT_RAM_35 = 256'h29BF2880288A1CC72980288A1CC702802880288A1CC72980288B1CC700102880;
defparam sp_inst_25.INIT_RAM_36 = 256'h5C000020028028BF293F002A5C000020028028BF500029BF02BF2880288A1CC7;
defparam sp_inst_25.INIT_RAM_37 = 256'h29BF02BF28BF57C100150280001502800280283F00150280004028BF29BF002A;
defparam sp_inst_25.INIT_RAM_38 = 256'h0010004002B11CC702BF28BF500029BF02805C0102802A0002951CC767FF28BF;
defparam sp_inst_25.INIT_RAM_39 = 256'h1CC7288028861CC763FF28BF29BF02BF28BF29800010004028BF02B01CC72880;
defparam sp_inst_25.INIT_RAM_3A = 256'h0340500029BF03BF140057E5028057B2298028851CC7298028861CC7298002AF;
defparam sp_inst_25.INIT_RAM_3B = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_3C = 256'h28BF034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_25.INIT_RAM_3D = 256'h5C0002802A00028F1CC72900028002AC1CC72900028002AD1CC747FF29BF02BF;
defparam sp_inst_25.INIT_RAM_3E = 256'h0015028002AE1C0002800280004028BF500029BF298028811CC7298028821CC7;
defparam sp_inst_25.INIT_RAM_3F = 256'h29BF0280298002BF4C00028028802880034067FF028028BF29BF028028BF57B8;

SP sp_inst_26 (
    .DO({sp_inst_26_dout_w[15:0],sp_inst_26_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_10}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_26.READ_MODE = 1'b0;
defparam sp_inst_26.WRITE_MODE = 2'b00;
defparam sp_inst_26.BIT_WIDTH = 16;
defparam sp_inst_26.BLK_SEL = 3'b001;
defparam sp_inst_26.RESET_MODE = "SYNC";
defparam sp_inst_26.INIT_RAM_00 = 256'h29BF03BF14006FFF028028BF29BF028028BF29800010004028BF02A91CC75000;
defparam sp_inst_26.INIT_RAM_01 = 256'h0340034003400340034003400340034003400340034003400340034003405000;
defparam sp_inst_26.INIT_RAM_02 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_26.INIT_RAM_03 = 256'h0280288003402900028002A61CC72900028002A71CC747FF29BF02BF28BF0340;
defparam sp_inst_26.INIT_RAM_04 = 256'h034057700380157F0280577202AA1C00028002B11C0002802980298002BF4C00;
defparam sp_inst_26.INIT_RAM_05 = 256'h157F0280577202A91C00028002B01C0002802980298002BF4C00028028802880;
defparam sp_inst_26.INIT_RAM_06 = 256'h02A81C00028002B01C0002802980298002BF4C000280288028800340576F0380;
defparam sp_inst_26.INIT_RAM_07 = 256'h02AF1C0002802980298002BF4C000280288028800340576F0380157F02805771;
defparam sp_inst_26.INIT_RAM_08 = 256'h2980298002BF4C000280288028800340576F0380157F0280577102A61C000280;
defparam sp_inst_26.INIT_RAM_09 = 256'h4C000280288028800340576F0380157F0280577102A51C00028002AE1C000280;
defparam sp_inst_26.INIT_RAM_0A = 256'h28800340576E0380157F0280577102A41C00028002AD1C0002802980298002BF;
defparam sp_inst_26.INIT_RAM_0B = 256'h0380157F0281577002A31C00028002AC1C0002802980298002BF4C0002802880;
defparam sp_inst_26.INIT_RAM_0C = 256'h577002A21C00028002AB1C0002802980298002BF4C000280288028800340576E;
defparam sp_inst_26.INIT_RAM_0D = 256'h028002AB1C0002802980298002BF4C000280288028800340576E0380157F0282;
defparam sp_inst_26.INIT_RAM_0E = 256'h02802980298002BF4C000280288028800340576D0380157F0284577002A01C00;
defparam sp_inst_26.INIT_RAM_0F = 256'h02BF4C000280288028800340576D0380157F0288576F029F1C00028102AA1C00;
defparam sp_inst_26.INIT_RAM_10 = 256'h288028800340576D0380157F0290576F029E1C00028102A91C00028029802980;
defparam sp_inst_26.INIT_RAM_11 = 256'h576C0380157F03A0576F029D1C00028102A81C0002802980298002BF4C000280;
defparam sp_inst_26.INIT_RAM_12 = 256'h1400576E029C1C00028102A71C0002802980298002BF4C000280288028800340;
defparam sp_inst_26.INIT_RAM_13 = 256'h1C00028102A71C0002802980298002BF4C000280288028800340576C0380157F;
defparam sp_inst_26.INIT_RAM_14 = 256'h1C0002802980298002BF4C000280288028800340576C0380157F1400576E029B;
defparam sp_inst_26.INIT_RAM_15 = 256'h298002BF4C000280288028800340576C0380157F1400576E02991C00028102A6;
defparam sp_inst_26.INIT_RAM_16 = 256'h0280288028800340576B0380157F1400576E02981C00028102A51C0002802980;
defparam sp_inst_26.INIT_RAM_17 = 256'h0340576B0380157F1400576D02971C00028102A41C0002802980298002BF4C00;
defparam sp_inst_26.INIT_RAM_18 = 256'h157F1400576D02961C00028102A31C0002802980298002BF4C00028028802880;
defparam sp_inst_26.INIT_RAM_19 = 256'h02951C00028102A31C0002802980298002BF4C000280288028800340576B0380;
defparam sp_inst_26.INIT_RAM_1A = 256'h02A21C0002802980298002BF4C000280288028800340576A0380157F1400576D;
defparam sp_inst_26.INIT_RAM_1B = 256'h2980298002BF4C000280288028800340576A0380157F1400576C02931C000281;
defparam sp_inst_26.INIT_RAM_1C = 256'h4C000280288028800340576A0380157F1400576C02921C00028202A11C000280;
defparam sp_inst_26.INIT_RAM_1D = 256'h2880034057690380157F1400576C02911C00028202A01C0002802980298002BF;
defparam sp_inst_26.INIT_RAM_1E = 256'h0380157F1400576C02901C000282029F1C0002802980298002BF4C0002802880;
defparam sp_inst_26.INIT_RAM_1F = 256'h576B028F1C000282029E1C0002802980298002BF4C0002802880288003405769;
defparam sp_inst_26.INIT_RAM_20 = 256'h0282029E1C0002802980298002BF4C00028028802880034057690380157F1401;
defparam sp_inst_26.INIT_RAM_21 = 256'h02802980298002BF4C00028028802880034057690380157F1402576B028D1C00;
defparam sp_inst_26.INIT_RAM_22 = 256'h02BF4C00028028802880034057680380157F1404576B028C1C000282029D1C00;
defparam sp_inst_26.INIT_RAM_23 = 256'h28802880034057680380157F1408576A028B1C000282029C1C00028029802980;
defparam sp_inst_26.INIT_RAM_24 = 256'h57680380157F1410576A028A1C000282029B1C0002802980298002BF4C000280;
defparam sp_inst_26.INIT_RAM_25 = 256'h1420576A02891C000282029A1C0002802980298002BF4C000280288028800340;
defparam sp_inst_26.INIT_RAM_26 = 256'h1C000282029A1C0002802980298002BF4C00028028802880034057670380157F;
defparam sp_inst_26.INIT_RAM_27 = 256'h1C0002802980298002BF4C00028028802880034057670380157F144057690288;
defparam sp_inst_26.INIT_RAM_28 = 256'h298002BF4C00028028802880034057670380157F1480576902861C0002820299;
defparam sp_inst_26.INIT_RAM_29 = 256'h028028802880034057670380157F1500576902851C00028302981C0002802980;
defparam sp_inst_26.INIT_RAM_2A = 256'h157F576802841C00028302971C00298014020380157F02802980298002BF4C00;
defparam sp_inst_26.INIT_RAM_2B = 256'h28BF28BF500029BF034029BF001428BF28BF29BF28800380157F29BF28800380;
defparam sp_inst_26.INIT_RAM_2C = 256'h6FFF028028BF29BF028028BF4C0028800010004028BF02861C00400003400017;
defparam sp_inst_26.INIT_RAM_2D = 256'h28800380157F298014000380157F02802980298002BF4C000280288028800340;
defparam sp_inst_26.INIT_RAM_2E = 256'h006F004428800380157F02802980298002BF4C000280288028800340576C29BF;
defparam sp_inst_26.INIT_RAM_2F = 256'h298002800380157F298014000380157F293F0340006728800380157F297F037F;
defparam sp_inst_26.INIT_RAM_30 = 256'h14000380157F0280298002BF4C000280288028800340576702BF1C0000152A7F;
defparam sp_inst_26.INIT_RAM_31 = 256'h28800380157F02802980298002BF4C00028028800340293F2A000380157F2980;
defparam sp_inst_26.INIT_RAM_32 = 256'h004028BF6800028028BF2980001414010380157F28800380157F29BF03400044;
defparam sp_inst_26.INIT_RAM_33 = 256'h157F576602BD1C00500029800380157F576602BD1C004C002880001002811C00;
defparam sp_inst_26.INIT_RAM_34 = 256'h02BF4C000280288028800340034050002980001403BF15FF0380157F28800380;
defparam sp_inst_26.INIT_RAM_35 = 256'h57A702844000001557A60284400003402A3F293F2A000380157F028029802980;
defparam sp_inst_26.INIT_RAM_36 = 256'h290002800380157F577100152A3F293F2880157F400003402A3F576602BB1C00;
defparam sp_inst_26.INIT_RAM_37 = 256'h02BF0380157F290002800380157F577100152A3F293F2880157F400003402A3F;
defparam sp_inst_26.INIT_RAM_38 = 256'h03405762576502B91C00576302802980298002BF4C0002802880288003402900;
defparam sp_inst_26.INIT_RAM_39 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C004C00028028802880;
defparam sp_inst_26.INIT_RAM_3A = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_26.INIT_RAM_3B = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_26.INIT_RAM_3C = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_26.INIT_RAM_3D = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_26.INIT_RAM_3E = 256'hB4D5BDFCBEFD0000202020204F2020201C001C001C001C001C001C001C001C00;
defparam sp_inst_26.INIT_RAM_3F = 256'h20ADCCF2B8ABCEB80000DCB0F1CFC6CEEBC80000B8D6D0D3CFC9D0B8000020F3;

SP sp_inst_27 (
    .DO({sp_inst_27_dout_w[15:0],sp_inst_27_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_11}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_27.READ_MODE = 1'b0;
defparam sp_inst_27.WRITE_MODE = 2'b00;
defparam sp_inst_27.BIT_WIDTH = 16;
defparam sp_inst_27.BLK_SEL = 3'b001;
defparam sp_inst_27.RESET_MODE = "SYNC";
defparam sp_inst_27.INIT_RAM_00 = 256'h000020D9CCE3D5D8CEB800002020ABCCBCCDB8D6000020FDCCF2CAABCEB80000;
defparam sp_inst_27.INIT_RAM_01 = 256'hB7D6000020DCCAA2BAF7CC20000020C6D6BDCBD1D3BB00002020E4C5BBB2B8D6;
defparam sp_inst_27.INIT_RAM_02 = 256'hDAC4E5B3000020DCCAE2CEB8BFE500002020A7CAA3C4BEC90000A7CEF6B3C5BA;
defparam sp_inst_27.INIT_RAM_03 = 256'hF7C6C4BCDECE00002020CEEDD2A8CE2000002020F6B3414CD0C10000BCCDD0D3;
defparam sp_inst_27.INIT_RAM_04 = 256'h2020FAC2C6CE2020000020F3B4EBD2BECAC7000020F3B4DDC4F7B4C400002020;
defparam sp_inst_27.INIT_RAM_05 = 256'h1C001C001C001C00003A000020F3D3EBC8B7BBB500002020F3CEB7D620200000;
defparam sp_inst_27.INIT_RAM_06 = 256'h001C0000221C000000005549231362007F2A147F140000070000000000001C00;
defparam sp_inst_27.INIT_RAM_07 = 256'h1214314B2100516100400000495102042000606008080800A000080808003E08;
defparam sp_inst_27.INIT_RAM_08 = 256'h020022411414140022140000000036361E290600494903050100494A39452700;
defparam sp_inst_27.INIT_RAM_09 = 256'h0041000008087A493E00090941497F00414122413E0049497C127C0059490609;
defparam sp_inst_27.INIT_RAM_0A = 256'h7F013149460019095E213E0009093E413E0008047F027F00404041227F004140;
defparam sp_inst_27.INIT_RAM_0B = 256'h40000102007F0000552A0041000049510708070008143F403F0040203F403F00;
defparam sp_inst_27.INIT_RAM_0C = 256'h0040000004087CA41800097E1854380044442044380044487854200002014040;
defparam sp_inst_27.INIT_RAM_0D = 256'h443F205448000408FC181800242438443800040878047C007F4100447F008480;
defparam sp_inst_27.INIT_RAM_0E = 256'hF80000000000000000001414141454647CA01C0010283C403C0040207C203C00;
defparam sp_inst_27.INIT_RAM_0F = 256'h00F00000FF200000FC880004040400404078000000000006060C000033000000;
defparam sp_inst_27.INIT_RAM_10 = 256'h1804004007000002E000000000000000000E1021242300008808001E031C0000;
defparam sp_inst_27.INIT_RAM_11 = 256'h0000000000700000000000011F010000F00000020F010040F080000018200000;
defparam sp_inst_27.INIT_RAM_12 = 256'hF810000F201000E0081000000618041800000000003000000000010101010000;
defparam sp_inst_27.INIT_RAM_13 = 256'h880800242404000020C0000E202000308808003024280070080800003F200000;
defparam sp_inst_27.INIT_RAM_14 = 256'h0810001C21220070088800003F0000080808000E201100008810000E20210008;
defparam sp_inst_27.INIT_RAM_15 = 256'h404000200402000840800000608000008000000030000000C000000F223100E0;
defparam sp_inst_27.INIT_RAM_16 = 256'h38C0000B242700E028C80000300000F008480001081000002010000404040040;
defparam sp_inst_27.INIT_RAM_17 = 256'h8888000F202000E008080008202000380808000E202000008888203802230000;
defparam sp_inst_27.INIT_RAM_18 = 256'hF808203F012108F8000800022020000008080000002000108888001820200010;
defparam sp_inst_27.INIT_RAM_19 = 256'h00F80030202000000008002001200008C088000080800008080800003F200000;
defparam sp_inst_27.INIT_RAM_1A = 256'h08080000012100F00808000F202000E00808003F002008F8C03000203F000008;
defparam sp_inst_27.INIT_RAM_1B = 256'h000800003F200018F808001C2120003808882030002000708888004F242400E0;
defparam sp_inst_27.INIT_RAM_1C = 256'h00C82030032C081880680003000700F8F8000000380708380088001F202008F8;
defparam sp_inst_27.INIT_RAM_1D = 256'h020200C001000000C03000407F000002FE00001821260008080800003F200008;
defparam sp_inst_27.INIT_RAM_1E = 256'h8080000000000000040280808080000000000000000000040204000040400000;
defparam sp_inst_27.INIT_RAM_1F = 256'h8080203F201100F880000011201100008000000E201100008000203F22240000;
defparam sp_inst_27.INIT_RAM_20 = 256'h9898203F002100008000006094940080808000003F201888F080001322220000;
defparam sp_inst_27.INIT_RAM_21 = 256'h808000003F200000F8080020022400800000000080800000800000003F200000;
defparam sp_inst_27.INIT_RAM_22 = 256'h8000000E20A100008000001F202000008080203F0021000080003F0000200080;
defparam sp_inst_27.INIT_RAM_23 = 256'h000000001F000000E08000192424008080800001213F0080008080FF20110080;
defparam sp_inst_27.INIT_RAM_24 = 256'h008000202E3100800080000F030C808080000001300E80800080203F20200080;
defparam sp_inst_27.INIT_RAM_25 = 256'h7C020000000000000000404000000202000000302C30008080800001708E8080;
defparam sp_inst_27.INIT_RAM_26 = 256'h000000000000000000000000000000000000000000000404010100003F400000;
defparam sp_inst_27.INIT_RAM_27 = 256'h000000000000000080C0C0C00000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_28 = 256'h0000000000000000000000000000FF0701000307000000000000000000000000;
defparam sp_inst_27.INIT_RAM_29 = 256'hFFFF3F1F00000000000000000000000000000000FFFFFF9F0F9FFFFFFE000000;
defparam sp_inst_27.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000071F7FFFF8F8;
defparam sp_inst_27.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2C = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_27.INIT_RAM_2D = 256'h1C001C001C001C001C001C001C00000000000000000000001C001C001C001C00;
defparam sp_inst_27.INIT_RAM_2E = 256'h3C201C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_27.INIT_RAM_2F = 256'h2E2E2E2E2E2E2E2E495F4F532E2E2E2E2E2E00000A0D20203A636620203A696C;
defparam sp_inst_27.INIT_RAM_30 = 256'h2E2E2E2E414641422E2E2E2E2E2E000078253A6C6E617965746E63752D2D0000;
defparam sp_inst_27.INIT_RAM_31 = 256'h656D20737265697200000A2E2E2E2E2E2E2E44412E2E2E2E2E2E00002E2E2E2E;
defparam sp_inst_27.INIT_RAM_32 = 256'h1C001C0000002E2E7572746E726163206D69657200000A2E7075657420726C63;
defparam sp_inst_27.INIT_RAM_33 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_27.INIT_RAM_34 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_27.INIT_RAM_35 = 256'h69741C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_27.INIT_RAM_36 = 256'h646E5F715F32697069740072646E5F715F31697069740072646E5F715F306970;
defparam sp_inst_27.INIT_RAM_37 = 256'h5F35697069740072646E5F715F34697069740072646E5F715F33697069740072;
defparam sp_inst_27.INIT_RAM_38 = 256'h69740072646E5F715F37697069740072646E5F715F36697069740072646E5F71;
defparam sp_inst_27.INIT_RAM_39 = 256'h646E5F715F32697069740072646E5F715F31697069740072646E5F715F306970;
defparam sp_inst_27.INIT_RAM_3A = 256'h5F35697069740072646E5F715F34697069740072646E5F715F33697069740072;
defparam sp_inst_27.INIT_RAM_3B = 256'h69740072646E5F715F37697069740072646E5F715F36697069740072646E5F71;
defparam sp_inst_27.INIT_RAM_3C = 256'h646E5F715F32697069740072646E5F715F31697069740072646E5F715F306970;
defparam sp_inst_27.INIT_RAM_3D = 256'h5F35697069740072646E5F715F34697069740072646E5F715F33697069740072;
defparam sp_inst_27.INIT_RAM_3E = 256'h69740072646E5F715F37697069740072646E5F715F36697069740072646E5F71;
defparam sp_inst_27.INIT_RAM_3F = 256'h646E5F715F32697069740072646E5F715F31697069740072646E5F715F306970;

SP sp_inst_28 (
    .DO({sp_inst_28_dout_w[15:0],sp_inst_28_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_12}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_28.READ_MODE = 1'b0;
defparam sp_inst_28.WRITE_MODE = 2'b00;
defparam sp_inst_28.BIT_WIDTH = 16;
defparam sp_inst_28.BLK_SEL = 3'b001;
defparam sp_inst_28.RESET_MODE = "SYNC";
defparam sp_inst_28.INIT_RAM_00 = 256'h5F35697069740072646E5F715F34697069740072646E5F715F33697069740072;
defparam sp_inst_28.INIT_RAM_01 = 256'h5F740072646E5F715F37697069740072646E5F715F36697069740072646E5F71;
defparam sp_inst_28.INIT_RAM_02 = 256'h1052325301E8000000001307FFFF80008000800080008000800000000072646E;
defparam sp_inst_28.INIT_RAM_03 = 256'h0202060100E08888007F121200E0888818CC494A0000FF494949FF0000004242;
defparam sp_inst_28.INIT_RAM_04 = 256'h62A2322200082909798929490040147F00241424000040000000000000000202;
defparam sp_inst_28.INIT_RAM_05 = 256'h44FF404000713F00304012220088888EC88863AC0000120A7E82132200008109;
defparam sp_inst_28.INIT_RAM_06 = 256'hE200E72C0008FF0900FF091F0000D20E00E027EC0000080400FF000000404444;
defparam sp_inst_28.INIT_RAM_07 = 256'h02005CE4000043427E42417A000C8414A69504440080100F4F807F01000020BF;
defparam sp_inst_28.INIT_RAM_08 = 256'hE200E72C0008FF0900FF091F0000D20E00E027EC003F48080800107F00808282;
defparam sp_inst_28.INIT_RAM_09 = 256'h7D55D5150080462843403F0000209E829EA0CC420080100F4F807F01000020BF;
defparam sp_inst_28.INIT_RAM_0A = 256'hC84ECC420000955515FF207F00405454545400CC00407F5555557F400000D555;
defparam sp_inst_28.INIT_RAM_0B = 256'h00E027EC000012121212017F00804A524A8610FF0040504F434C1F20000048C8;
defparam sp_inst_28.INIT_RAM_0C = 256'h8E8908080080100F4F807F01000020BFE200E72C0008FF0900FF091F0000D20E;
defparam sp_inst_28.INIT_RAM_0D = 256'h545400CC00F8100C10102060001010101090909000003F400000204000088888;
defparam sp_inst_28.INIT_RAM_0E = 256'h1CE2000000005F0012FFFF090010941254C8C81F0000955515FF207F00405454;
defparam sp_inst_28.INIT_RAM_0F = 256'h02005CE4000043427E42417A000C8414A69504440080300C0000102000000000;
defparam sp_inst_28.INIT_RAM_10 = 256'hE200E72C0008FF0900FF091F0000D20E00E027EC003F48080800107F00808282;
defparam sp_inst_28.INIT_RAM_11 = 256'h2040FA02008121110103214100001010FF101E300080100F4F807F01000020BF;
defparam sp_inst_28.INIT_RAM_12 = 256'h1008F80800F81816801F001F00080908088888F80080160840800F3000101010;
defparam sp_inst_28.INIT_RAM_13 = 256'hFE2222FE00804141294500FF00042424242407F80000804030481F1000001010;
defparam sp_inst_28.INIT_RAM_14 = 256'hFE00FC840000F84B4A4AFF00006226A2BAA2A223000082427F02021F00002222;
defparam sp_inst_28.INIT_RAM_15 = 256'h49FFCC42000020200E10408F00005E5252525EC00040447F44401F20000092FE;
defparam sp_inst_28.INIT_RAM_16 = 256'h24FCCC42000040407F40404000004040FF40407C00404241485F1F2000004949;
defparam sp_inst_28.INIT_RAM_17 = 256'h30408444000020202424207F00000202121202FE0040454250471F2000002222;
defparam sp_inst_28.INIT_RAM_18 = 256'h7F4044420040427F444F1F20000004FC04FCCC42008018061820010600000808;
defparam sp_inst_28.INIT_RAM_19 = 256'h24FCCC420000213F7F0000000008086818200000007840400000204000404850;
defparam sp_inst_28.INIT_RAM_1A = 256'h52928C02000020202424207F00000202121202FE0040454250471F2000002222;
defparam sp_inst_28.INIT_RAM_1B = 256'h3D6424FC00002020007F0F300000080800F0FF10003130084018017E00105232;
defparam sp_inst_28.INIT_RAM_1C = 256'h28105A220000955515FF017E0040545454548C02001012121212100F00042424;
defparam sp_inst_28.INIT_RAM_1D = 256'h49497F00000040404040403F0000FE82828282E200000501410D080400202824;
defparam sp_inst_28.INIT_RAM_1E = 256'h3F00FF100001FC444544FC0000004222FA12828200818989FF811D2100007F49;
defparam sp_inst_28.INIT_RAM_1F = 256'h545400CC00802116214012220000F808F80863AC00004949FF007F8200704444;
defparam sp_inst_28.INIT_RAM_20 = 256'hFC2424240000281084807F810098888E8898FF100000955515FF207F00405454;
defparam sp_inst_28.INIT_RAM_21 = 256'h9292928200004949FF007F82007044443F00FF10000202027F82020200002322;
defparam sp_inst_28.INIT_RAM_22 = 256'h3F00FF100080300C00001020000000001CE20000004024187F8024220080FE92;
defparam sp_inst_28.INIT_RAM_23 = 256'h088888F800802116214012220000F808F80863AC00004949FF007F8200704444;
defparam sp_inst_28.INIT_RAM_24 = 256'hFF101E300000804030481F10000010101008F80800F81816801F001F00080908;
defparam sp_inst_28.INIT_RAM_25 = 256'h9292927E0080160840800F30001010102040FA02008121110103214100001010;
defparam sp_inst_28.INIT_RAM_26 = 256'h545400CC00002212FF02023E0018EAACAFA8EA08000808FE0808284800009E92;
defparam sp_inst_28.INIT_RAM_27 = 256'h2424FC0000004909FF00FF010000203FE200FEA40000955515FF207F00405454;
defparam sp_inst_28.INIT_RAM_28 = 256'h9090CC4200048444070404FF00029292FE9292F2000042424242071800202322;
defparam sp_inst_28.INIT_RAM_29 = 256'h5455FC0000000404FF04040F00001010FF1010F000F00E013F603F00001010FF;
defparam sp_inst_28.INIT_RAM_2A = 256'h20408282000080403040FF0000808780B040F86000007F82121223420040FC54;
defparam sp_inst_28.INIT_RAM_2B = 256'h000000000040417F7F403F00000404FCC404CC420040604E4440844800404C43;
defparam sp_inst_28.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_29 (
    .DO({sp_inst_29_dout_w[15:0],sp_inst_29_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_13}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_29.READ_MODE = 1'b0;
defparam sp_inst_29.WRITE_MODE = 2'b00;
defparam sp_inst_29.BIT_WIDTH = 16;
defparam sp_inst_29.BLK_SEL = 3'b001;
defparam sp_inst_29.RESET_MODE = "SYNC";
defparam sp_inst_29.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_30 (
    .DO({sp_inst_30_dout_w[15:0],sp_inst_30_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_14}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_30.READ_MODE = 1'b0;
defparam sp_inst_30.WRITE_MODE = 2'b00;
defparam sp_inst_30.BIT_WIDTH = 16;
defparam sp_inst_30.BLK_SEL = 3'b001;
defparam sp_inst_30.RESET_MODE = "SYNC";
defparam sp_inst_30.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_31 (
    .DO({sp_inst_31_dout_w[15:0],sp_inst_31_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_15}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_31.READ_MODE = 1'b0;
defparam sp_inst_31.WRITE_MODE = 2'b00;
defparam sp_inst_31.BIT_WIDTH = 16;
defparam sp_inst_31.BLK_SEL = 3'b001;
defparam sp_inst_31.RESET_MODE = "SYNC";
defparam sp_inst_31.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_3 (
  .Q(dff_q_3),
  .D(ad[10]),
  .CLK(clk),
  .CE(ce_w),
  .RESET(gw_gnd)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(sp_inst_0_dout[0]),
  .I1(sp_inst_1_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(sp_inst_2_dout[0]),
  .I1(sp_inst_3_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(sp_inst_4_dout[0]),
  .I1(sp_inst_5_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(sp_inst_6_dout[0]),
  .I1(sp_inst_7_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(sp_inst_8_dout[0]),
  .I1(sp_inst_9_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(sp_inst_10_dout[0]),
  .I1(sp_inst_11_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(sp_inst_12_dout[0]),
  .I1(sp_inst_13_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(sp_inst_14_dout[0]),
  .I1(sp_inst_15_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_2)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_2)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_2)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(dff_q_2)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(dff_q_1)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_1)
);
MUX2 mux_inst_14 (
  .O(dout[0]),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_0)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(sp_inst_0_dout[1]),
  .I1(sp_inst_1_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(sp_inst_2_dout[1]),
  .I1(sp_inst_3_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(sp_inst_4_dout[1]),
  .I1(sp_inst_5_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(sp_inst_6_dout[1]),
  .I1(sp_inst_7_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(sp_inst_8_dout[1]),
  .I1(sp_inst_9_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(sp_inst_10_dout[1]),
  .I1(sp_inst_11_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(sp_inst_12_dout[1]),
  .I1(sp_inst_13_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(sp_inst_14_dout[1]),
  .I1(sp_inst_15_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(mux_o_15),
  .I1(mux_o_16),
  .S0(dff_q_2)
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(mux_o_17),
  .I1(mux_o_18),
  .S0(dff_q_2)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(mux_o_19),
  .I1(mux_o_20),
  .S0(dff_q_2)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(mux_o_21),
  .I1(mux_o_22),
  .S0(dff_q_2)
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(mux_o_23),
  .I1(mux_o_24),
  .S0(dff_q_1)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(mux_o_25),
  .I1(mux_o_26),
  .S0(dff_q_1)
);
MUX2 mux_inst_29 (
  .O(dout[1]),
  .I0(mux_o_27),
  .I1(mux_o_28),
  .S0(dff_q_0)
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(sp_inst_0_dout[2]),
  .I1(sp_inst_1_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(sp_inst_2_dout[2]),
  .I1(sp_inst_3_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(sp_inst_4_dout[2]),
  .I1(sp_inst_5_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(sp_inst_6_dout[2]),
  .I1(sp_inst_7_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(sp_inst_8_dout[2]),
  .I1(sp_inst_9_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(sp_inst_10_dout[2]),
  .I1(sp_inst_11_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(sp_inst_12_dout[2]),
  .I1(sp_inst_13_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(sp_inst_14_dout[2]),
  .I1(sp_inst_15_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(dff_q_2)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(dff_q_2)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_34),
  .I1(mux_o_35),
  .S0(dff_q_2)
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(mux_o_36),
  .I1(mux_o_37),
  .S0(dff_q_2)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(dff_q_1)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(dff_q_1)
);
MUX2 mux_inst_44 (
  .O(dout[2]),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(dff_q_0)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(sp_inst_0_dout[3]),
  .I1(sp_inst_1_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(sp_inst_2_dout[3]),
  .I1(sp_inst_3_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(sp_inst_4_dout[3]),
  .I1(sp_inst_5_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(sp_inst_6_dout[3]),
  .I1(sp_inst_7_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(sp_inst_8_dout[3]),
  .I1(sp_inst_9_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(sp_inst_10_dout[3]),
  .I1(sp_inst_11_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(sp_inst_12_dout[3]),
  .I1(sp_inst_13_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(sp_inst_14_dout[3]),
  .I1(sp_inst_15_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(dff_q_2)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_47),
  .I1(mux_o_48),
  .S0(dff_q_2)
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(dff_q_2)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(mux_o_51),
  .I1(mux_o_52),
  .S0(dff_q_2)
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(mux_o_53),
  .I1(mux_o_54),
  .S0(dff_q_1)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(mux_o_55),
  .I1(mux_o_56),
  .S0(dff_q_1)
);
MUX2 mux_inst_59 (
  .O(dout[3]),
  .I0(mux_o_57),
  .I1(mux_o_58),
  .S0(dff_q_0)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(sp_inst_0_dout[4]),
  .I1(sp_inst_1_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(sp_inst_2_dout[4]),
  .I1(sp_inst_3_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(sp_inst_4_dout[4]),
  .I1(sp_inst_5_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(sp_inst_6_dout[4]),
  .I1(sp_inst_7_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(sp_inst_8_dout[4]),
  .I1(sp_inst_9_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(sp_inst_10_dout[4]),
  .I1(sp_inst_11_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(sp_inst_12_dout[4]),
  .I1(sp_inst_13_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(sp_inst_14_dout[4]),
  .I1(sp_inst_15_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(dff_q_2)
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(dff_q_2)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(mux_o_64),
  .I1(mux_o_65),
  .S0(dff_q_2)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(dff_q_2)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(mux_o_68),
  .I1(mux_o_69),
  .S0(dff_q_1)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(dff_q_1)
);
MUX2 mux_inst_74 (
  .O(dout[4]),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(dff_q_0)
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(sp_inst_0_dout[5]),
  .I1(sp_inst_1_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(sp_inst_2_dout[5]),
  .I1(sp_inst_3_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(sp_inst_4_dout[5]),
  .I1(sp_inst_5_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(sp_inst_6_dout[5]),
  .I1(sp_inst_7_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(sp_inst_8_dout[5]),
  .I1(sp_inst_9_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(sp_inst_10_dout[5]),
  .I1(sp_inst_11_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(sp_inst_12_dout[5]),
  .I1(sp_inst_13_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(sp_inst_14_dout[5]),
  .I1(sp_inst_15_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(mux_o_75),
  .I1(mux_o_76),
  .S0(dff_q_2)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(dff_q_2)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(dff_q_2)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(dff_q_2)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(mux_o_83),
  .I1(mux_o_84),
  .S0(dff_q_1)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(dff_q_1)
);
MUX2 mux_inst_89 (
  .O(dout[5]),
  .I0(mux_o_87),
  .I1(mux_o_88),
  .S0(dff_q_0)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(sp_inst_0_dout[6]),
  .I1(sp_inst_1_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(sp_inst_2_dout[6]),
  .I1(sp_inst_3_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(sp_inst_4_dout[6]),
  .I1(sp_inst_5_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(sp_inst_6_dout[6]),
  .I1(sp_inst_7_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(sp_inst_8_dout[6]),
  .I1(sp_inst_9_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(sp_inst_10_dout[6]),
  .I1(sp_inst_11_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(sp_inst_12_dout[6]),
  .I1(sp_inst_13_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(sp_inst_14_dout[6]),
  .I1(sp_inst_15_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(dff_q_2)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(dff_q_2)
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(mux_o_94),
  .I1(mux_o_95),
  .S0(dff_q_2)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_96),
  .I1(mux_o_97),
  .S0(dff_q_2)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_98),
  .I1(mux_o_99),
  .S0(dff_q_1)
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(mux_o_100),
  .I1(mux_o_101),
  .S0(dff_q_1)
);
MUX2 mux_inst_104 (
  .O(dout[6]),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(dff_q_0)
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(sp_inst_0_dout[7]),
  .I1(sp_inst_1_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(sp_inst_2_dout[7]),
  .I1(sp_inst_3_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(sp_inst_4_dout[7]),
  .I1(sp_inst_5_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(sp_inst_6_dout[7]),
  .I1(sp_inst_7_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(sp_inst_8_dout[7]),
  .I1(sp_inst_9_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(sp_inst_10_dout[7]),
  .I1(sp_inst_11_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(sp_inst_12_dout[7]),
  .I1(sp_inst_13_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(sp_inst_14_dout[7]),
  .I1(sp_inst_15_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(dff_q_2)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(dff_q_2)
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(dff_q_2)
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_111),
  .I1(mux_o_112),
  .S0(dff_q_2)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_113),
  .I1(mux_o_114),
  .S0(dff_q_1)
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_115),
  .I1(mux_o_116),
  .S0(dff_q_1)
);
MUX2 mux_inst_119 (
  .O(dout[7]),
  .I0(mux_o_117),
  .I1(mux_o_118),
  .S0(dff_q_0)
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(sp_inst_0_dout[8]),
  .I1(sp_inst_1_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(sp_inst_2_dout[8]),
  .I1(sp_inst_3_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(sp_inst_4_dout[8]),
  .I1(sp_inst_5_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(sp_inst_6_dout[8]),
  .I1(sp_inst_7_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(sp_inst_8_dout[8]),
  .I1(sp_inst_9_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_125 (
  .O(mux_o_125),
  .I0(sp_inst_10_dout[8]),
  .I1(sp_inst_11_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(sp_inst_12_dout[8]),
  .I1(sp_inst_13_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(sp_inst_14_dout[8]),
  .I1(sp_inst_15_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(mux_o_120),
  .I1(mux_o_121),
  .S0(dff_q_2)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(mux_o_122),
  .I1(mux_o_123),
  .S0(dff_q_2)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(mux_o_124),
  .I1(mux_o_125),
  .S0(dff_q_2)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(dff_q_2)
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(dff_q_1)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(dff_q_1)
);
MUX2 mux_inst_134 (
  .O(dout[8]),
  .I0(mux_o_132),
  .I1(mux_o_133),
  .S0(dff_q_0)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(sp_inst_0_dout[9]),
  .I1(sp_inst_1_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(sp_inst_2_dout[9]),
  .I1(sp_inst_3_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(sp_inst_4_dout[9]),
  .I1(sp_inst_5_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(sp_inst_6_dout[9]),
  .I1(sp_inst_7_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(sp_inst_8_dout[9]),
  .I1(sp_inst_9_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(sp_inst_10_dout[9]),
  .I1(sp_inst_11_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(sp_inst_12_dout[9]),
  .I1(sp_inst_13_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(sp_inst_14_dout[9]),
  .I1(sp_inst_15_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(mux_o_135),
  .I1(mux_o_136),
  .S0(dff_q_2)
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(dff_q_2)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(mux_o_139),
  .I1(mux_o_140),
  .S0(dff_q_2)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(mux_o_141),
  .I1(mux_o_142),
  .S0(dff_q_2)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(mux_o_143),
  .I1(mux_o_144),
  .S0(dff_q_1)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(mux_o_145),
  .I1(mux_o_146),
  .S0(dff_q_1)
);
MUX2 mux_inst_149 (
  .O(dout[9]),
  .I0(mux_o_147),
  .I1(mux_o_148),
  .S0(dff_q_0)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(sp_inst_0_dout[10]),
  .I1(sp_inst_1_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(sp_inst_2_dout[10]),
  .I1(sp_inst_3_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(sp_inst_4_dout[10]),
  .I1(sp_inst_5_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(sp_inst_6_dout[10]),
  .I1(sp_inst_7_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(sp_inst_8_dout[10]),
  .I1(sp_inst_9_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(sp_inst_10_dout[10]),
  .I1(sp_inst_11_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(sp_inst_12_dout[10]),
  .I1(sp_inst_13_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(sp_inst_14_dout[10]),
  .I1(sp_inst_15_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(mux_o_150),
  .I1(mux_o_151),
  .S0(dff_q_2)
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(mux_o_152),
  .I1(mux_o_153),
  .S0(dff_q_2)
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(mux_o_154),
  .I1(mux_o_155),
  .S0(dff_q_2)
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(mux_o_156),
  .I1(mux_o_157),
  .S0(dff_q_2)
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(mux_o_158),
  .I1(mux_o_159),
  .S0(dff_q_1)
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(mux_o_160),
  .I1(mux_o_161),
  .S0(dff_q_1)
);
MUX2 mux_inst_164 (
  .O(dout[10]),
  .I0(mux_o_162),
  .I1(mux_o_163),
  .S0(dff_q_0)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(sp_inst_0_dout[11]),
  .I1(sp_inst_1_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(sp_inst_2_dout[11]),
  .I1(sp_inst_3_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(sp_inst_4_dout[11]),
  .I1(sp_inst_5_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(sp_inst_6_dout[11]),
  .I1(sp_inst_7_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(sp_inst_8_dout[11]),
  .I1(sp_inst_9_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(sp_inst_10_dout[11]),
  .I1(sp_inst_11_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(sp_inst_12_dout[11]),
  .I1(sp_inst_13_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(sp_inst_14_dout[11]),
  .I1(sp_inst_15_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(dff_q_2)
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(mux_o_167),
  .I1(mux_o_168),
  .S0(dff_q_2)
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(mux_o_169),
  .I1(mux_o_170),
  .S0(dff_q_2)
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(mux_o_171),
  .I1(mux_o_172),
  .S0(dff_q_2)
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(mux_o_173),
  .I1(mux_o_174),
  .S0(dff_q_1)
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(mux_o_175),
  .I1(mux_o_176),
  .S0(dff_q_1)
);
MUX2 mux_inst_179 (
  .O(dout[11]),
  .I0(mux_o_177),
  .I1(mux_o_178),
  .S0(dff_q_0)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(sp_inst_0_dout[12]),
  .I1(sp_inst_1_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(sp_inst_2_dout[12]),
  .I1(sp_inst_3_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(sp_inst_4_dout[12]),
  .I1(sp_inst_5_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(sp_inst_6_dout[12]),
  .I1(sp_inst_7_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(sp_inst_8_dout[12]),
  .I1(sp_inst_9_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(sp_inst_10_dout[12]),
  .I1(sp_inst_11_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(sp_inst_12_dout[12]),
  .I1(sp_inst_13_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(sp_inst_14_dout[12]),
  .I1(sp_inst_15_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(mux_o_180),
  .I1(mux_o_181),
  .S0(dff_q_2)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(mux_o_182),
  .I1(mux_o_183),
  .S0(dff_q_2)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(mux_o_184),
  .I1(mux_o_185),
  .S0(dff_q_2)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(dff_q_2)
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(mux_o_188),
  .I1(mux_o_189),
  .S0(dff_q_1)
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(mux_o_190),
  .I1(mux_o_191),
  .S0(dff_q_1)
);
MUX2 mux_inst_194 (
  .O(dout[12]),
  .I0(mux_o_192),
  .I1(mux_o_193),
  .S0(dff_q_0)
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(sp_inst_0_dout[13]),
  .I1(sp_inst_1_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(sp_inst_2_dout[13]),
  .I1(sp_inst_3_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(sp_inst_4_dout[13]),
  .I1(sp_inst_5_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(sp_inst_6_dout[13]),
  .I1(sp_inst_7_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(sp_inst_8_dout[13]),
  .I1(sp_inst_9_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(sp_inst_10_dout[13]),
  .I1(sp_inst_11_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(sp_inst_12_dout[13]),
  .I1(sp_inst_13_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(sp_inst_14_dout[13]),
  .I1(sp_inst_15_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_195),
  .I1(mux_o_196),
  .S0(dff_q_2)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(mux_o_197),
  .I1(mux_o_198),
  .S0(dff_q_2)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_199),
  .I1(mux_o_200),
  .S0(dff_q_2)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_201),
  .I1(mux_o_202),
  .S0(dff_q_2)
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(mux_o_203),
  .I1(mux_o_204),
  .S0(dff_q_1)
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(dff_q_1)
);
MUX2 mux_inst_209 (
  .O(dout[13]),
  .I0(mux_o_207),
  .I1(mux_o_208),
  .S0(dff_q_0)
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(sp_inst_0_dout[14]),
  .I1(sp_inst_1_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(sp_inst_2_dout[14]),
  .I1(sp_inst_3_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(sp_inst_4_dout[14]),
  .I1(sp_inst_5_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(sp_inst_6_dout[14]),
  .I1(sp_inst_7_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(sp_inst_8_dout[14]),
  .I1(sp_inst_9_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(sp_inst_10_dout[14]),
  .I1(sp_inst_11_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(sp_inst_12_dout[14]),
  .I1(sp_inst_13_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(sp_inst_14_dout[14]),
  .I1(sp_inst_15_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(mux_o_210),
  .I1(mux_o_211),
  .S0(dff_q_2)
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(mux_o_212),
  .I1(mux_o_213),
  .S0(dff_q_2)
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(mux_o_214),
  .I1(mux_o_215),
  .S0(dff_q_2)
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(mux_o_216),
  .I1(mux_o_217),
  .S0(dff_q_2)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(mux_o_218),
  .I1(mux_o_219),
  .S0(dff_q_1)
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(mux_o_220),
  .I1(mux_o_221),
  .S0(dff_q_1)
);
MUX2 mux_inst_224 (
  .O(dout[14]),
  .I0(mux_o_222),
  .I1(mux_o_223),
  .S0(dff_q_0)
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(sp_inst_0_dout[15]),
  .I1(sp_inst_1_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(sp_inst_2_dout[15]),
  .I1(sp_inst_3_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(sp_inst_4_dout[15]),
  .I1(sp_inst_5_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(sp_inst_6_dout[15]),
  .I1(sp_inst_7_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(sp_inst_8_dout[15]),
  .I1(sp_inst_9_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(sp_inst_10_dout[15]),
  .I1(sp_inst_11_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(sp_inst_12_dout[15]),
  .I1(sp_inst_13_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(sp_inst_14_dout[15]),
  .I1(sp_inst_15_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_225),
  .I1(mux_o_226),
  .S0(dff_q_2)
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(mux_o_227),
  .I1(mux_o_228),
  .S0(dff_q_2)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_229),
  .I1(mux_o_230),
  .S0(dff_q_2)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(dff_q_2)
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(dff_q_1)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_1)
);
MUX2 mux_inst_239 (
  .O(dout[15]),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(dff_q_0)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(sp_inst_16_dout[16]),
  .I1(sp_inst_17_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(sp_inst_18_dout[16]),
  .I1(sp_inst_19_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(sp_inst_20_dout[16]),
  .I1(sp_inst_21_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(sp_inst_22_dout[16]),
  .I1(sp_inst_23_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(sp_inst_24_dout[16]),
  .I1(sp_inst_25_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(sp_inst_26_dout[16]),
  .I1(sp_inst_27_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(sp_inst_28_dout[16]),
  .I1(sp_inst_29_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(sp_inst_30_dout[16]),
  .I1(sp_inst_31_dout[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(mux_o_240),
  .I1(mux_o_241),
  .S0(dff_q_2)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_242),
  .I1(mux_o_243),
  .S0(dff_q_2)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_244),
  .I1(mux_o_245),
  .S0(dff_q_2)
);
MUX2 mux_inst_251 (
  .O(mux_o_251),
  .I0(mux_o_246),
  .I1(mux_o_247),
  .S0(dff_q_2)
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(mux_o_248),
  .I1(mux_o_249),
  .S0(dff_q_1)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(mux_o_250),
  .I1(mux_o_251),
  .S0(dff_q_1)
);
MUX2 mux_inst_254 (
  .O(dout[16]),
  .I0(mux_o_252),
  .I1(mux_o_253),
  .S0(dff_q_0)
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(sp_inst_16_dout[17]),
  .I1(sp_inst_17_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(sp_inst_18_dout[17]),
  .I1(sp_inst_19_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(sp_inst_20_dout[17]),
  .I1(sp_inst_21_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(sp_inst_22_dout[17]),
  .I1(sp_inst_23_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(sp_inst_24_dout[17]),
  .I1(sp_inst_25_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(sp_inst_26_dout[17]),
  .I1(sp_inst_27_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(sp_inst_28_dout[17]),
  .I1(sp_inst_29_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(sp_inst_30_dout[17]),
  .I1(sp_inst_31_dout[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(mux_o_255),
  .I1(mux_o_256),
  .S0(dff_q_2)
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(mux_o_257),
  .I1(mux_o_258),
  .S0(dff_q_2)
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(mux_o_259),
  .I1(mux_o_260),
  .S0(dff_q_2)
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(mux_o_261),
  .I1(mux_o_262),
  .S0(dff_q_2)
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(mux_o_263),
  .I1(mux_o_264),
  .S0(dff_q_1)
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(mux_o_265),
  .I1(mux_o_266),
  .S0(dff_q_1)
);
MUX2 mux_inst_269 (
  .O(dout[17]),
  .I0(mux_o_267),
  .I1(mux_o_268),
  .S0(dff_q_0)
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(sp_inst_16_dout[18]),
  .I1(sp_inst_17_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(sp_inst_18_dout[18]),
  .I1(sp_inst_19_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_272 (
  .O(mux_o_272),
  .I0(sp_inst_20_dout[18]),
  .I1(sp_inst_21_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(sp_inst_22_dout[18]),
  .I1(sp_inst_23_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(sp_inst_24_dout[18]),
  .I1(sp_inst_25_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(sp_inst_26_dout[18]),
  .I1(sp_inst_27_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(sp_inst_28_dout[18]),
  .I1(sp_inst_29_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(sp_inst_30_dout[18]),
  .I1(sp_inst_31_dout[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(dff_q_2)
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(mux_o_272),
  .I1(mux_o_273),
  .S0(dff_q_2)
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(mux_o_274),
  .I1(mux_o_275),
  .S0(dff_q_2)
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(mux_o_276),
  .I1(mux_o_277),
  .S0(dff_q_2)
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(mux_o_278),
  .I1(mux_o_279),
  .S0(dff_q_1)
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(mux_o_280),
  .I1(mux_o_281),
  .S0(dff_q_1)
);
MUX2 mux_inst_284 (
  .O(dout[18]),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(dff_q_0)
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(sp_inst_16_dout[19]),
  .I1(sp_inst_17_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(sp_inst_18_dout[19]),
  .I1(sp_inst_19_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(sp_inst_20_dout[19]),
  .I1(sp_inst_21_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(sp_inst_22_dout[19]),
  .I1(sp_inst_23_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(sp_inst_24_dout[19]),
  .I1(sp_inst_25_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(sp_inst_26_dout[19]),
  .I1(sp_inst_27_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(sp_inst_28_dout[19]),
  .I1(sp_inst_29_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(sp_inst_30_dout[19]),
  .I1(sp_inst_31_dout[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(mux_o_285),
  .I1(mux_o_286),
  .S0(dff_q_2)
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(mux_o_287),
  .I1(mux_o_288),
  .S0(dff_q_2)
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(mux_o_289),
  .I1(mux_o_290),
  .S0(dff_q_2)
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(mux_o_291),
  .I1(mux_o_292),
  .S0(dff_q_2)
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(mux_o_293),
  .I1(mux_o_294),
  .S0(dff_q_1)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(mux_o_295),
  .I1(mux_o_296),
  .S0(dff_q_1)
);
MUX2 mux_inst_299 (
  .O(dout[19]),
  .I0(mux_o_297),
  .I1(mux_o_298),
  .S0(dff_q_0)
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(sp_inst_16_dout[20]),
  .I1(sp_inst_17_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(sp_inst_18_dout[20]),
  .I1(sp_inst_19_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(sp_inst_20_dout[20]),
  .I1(sp_inst_21_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(sp_inst_22_dout[20]),
  .I1(sp_inst_23_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(sp_inst_24_dout[20]),
  .I1(sp_inst_25_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(sp_inst_26_dout[20]),
  .I1(sp_inst_27_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(sp_inst_28_dout[20]),
  .I1(sp_inst_29_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(sp_inst_30_dout[20]),
  .I1(sp_inst_31_dout[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(mux_o_300),
  .I1(mux_o_301),
  .S0(dff_q_2)
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(mux_o_302),
  .I1(mux_o_303),
  .S0(dff_q_2)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(mux_o_304),
  .I1(mux_o_305),
  .S0(dff_q_2)
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(mux_o_306),
  .I1(mux_o_307),
  .S0(dff_q_2)
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(mux_o_308),
  .I1(mux_o_309),
  .S0(dff_q_1)
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(dff_q_1)
);
MUX2 mux_inst_314 (
  .O(dout[20]),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(dff_q_0)
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(sp_inst_16_dout[21]),
  .I1(sp_inst_17_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(sp_inst_18_dout[21]),
  .I1(sp_inst_19_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(sp_inst_20_dout[21]),
  .I1(sp_inst_21_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(sp_inst_22_dout[21]),
  .I1(sp_inst_23_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(sp_inst_24_dout[21]),
  .I1(sp_inst_25_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(sp_inst_26_dout[21]),
  .I1(sp_inst_27_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(sp_inst_28_dout[21]),
  .I1(sp_inst_29_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(sp_inst_30_dout[21]),
  .I1(sp_inst_31_dout[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(mux_o_315),
  .I1(mux_o_316),
  .S0(dff_q_2)
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(mux_o_317),
  .I1(mux_o_318),
  .S0(dff_q_2)
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(mux_o_319),
  .I1(mux_o_320),
  .S0(dff_q_2)
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(mux_o_321),
  .I1(mux_o_322),
  .S0(dff_q_2)
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(mux_o_323),
  .I1(mux_o_324),
  .S0(dff_q_1)
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(mux_o_325),
  .I1(mux_o_326),
  .S0(dff_q_1)
);
MUX2 mux_inst_329 (
  .O(dout[21]),
  .I0(mux_o_327),
  .I1(mux_o_328),
  .S0(dff_q_0)
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(sp_inst_16_dout[22]),
  .I1(sp_inst_17_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(sp_inst_18_dout[22]),
  .I1(sp_inst_19_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(sp_inst_20_dout[22]),
  .I1(sp_inst_21_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(sp_inst_22_dout[22]),
  .I1(sp_inst_23_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(sp_inst_24_dout[22]),
  .I1(sp_inst_25_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(sp_inst_26_dout[22]),
  .I1(sp_inst_27_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(sp_inst_28_dout[22]),
  .I1(sp_inst_29_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(sp_inst_30_dout[22]),
  .I1(sp_inst_31_dout[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(mux_o_330),
  .I1(mux_o_331),
  .S0(dff_q_2)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(mux_o_332),
  .I1(mux_o_333),
  .S0(dff_q_2)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(mux_o_334),
  .I1(mux_o_335),
  .S0(dff_q_2)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(mux_o_336),
  .I1(mux_o_337),
  .S0(dff_q_2)
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(mux_o_338),
  .I1(mux_o_339),
  .S0(dff_q_1)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(mux_o_340),
  .I1(mux_o_341),
  .S0(dff_q_1)
);
MUX2 mux_inst_344 (
  .O(dout[22]),
  .I0(mux_o_342),
  .I1(mux_o_343),
  .S0(dff_q_0)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(sp_inst_16_dout[23]),
  .I1(sp_inst_17_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(sp_inst_18_dout[23]),
  .I1(sp_inst_19_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(sp_inst_20_dout[23]),
  .I1(sp_inst_21_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(sp_inst_22_dout[23]),
  .I1(sp_inst_23_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_349 (
  .O(mux_o_349),
  .I0(sp_inst_24_dout[23]),
  .I1(sp_inst_25_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(sp_inst_26_dout[23]),
  .I1(sp_inst_27_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(sp_inst_28_dout[23]),
  .I1(sp_inst_29_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(sp_inst_30_dout[23]),
  .I1(sp_inst_31_dout[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(mux_o_345),
  .I1(mux_o_346),
  .S0(dff_q_2)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(dff_q_2)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(mux_o_349),
  .I1(mux_o_350),
  .S0(dff_q_2)
);
MUX2 mux_inst_356 (
  .O(mux_o_356),
  .I0(mux_o_351),
  .I1(mux_o_352),
  .S0(dff_q_2)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_353),
  .I1(mux_o_354),
  .S0(dff_q_1)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_355),
  .I1(mux_o_356),
  .S0(dff_q_1)
);
MUX2 mux_inst_359 (
  .O(dout[23]),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(dff_q_0)
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(sp_inst_16_dout[24]),
  .I1(sp_inst_17_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(sp_inst_18_dout[24]),
  .I1(sp_inst_19_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(sp_inst_20_dout[24]),
  .I1(sp_inst_21_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_363 (
  .O(mux_o_363),
  .I0(sp_inst_22_dout[24]),
  .I1(sp_inst_23_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(sp_inst_24_dout[24]),
  .I1(sp_inst_25_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(sp_inst_26_dout[24]),
  .I1(sp_inst_27_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(sp_inst_28_dout[24]),
  .I1(sp_inst_29_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(sp_inst_30_dout[24]),
  .I1(sp_inst_31_dout[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(mux_o_360),
  .I1(mux_o_361),
  .S0(dff_q_2)
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(mux_o_362),
  .I1(mux_o_363),
  .S0(dff_q_2)
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(mux_o_364),
  .I1(mux_o_365),
  .S0(dff_q_2)
);
MUX2 mux_inst_371 (
  .O(mux_o_371),
  .I0(mux_o_366),
  .I1(mux_o_367),
  .S0(dff_q_2)
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(mux_o_368),
  .I1(mux_o_369),
  .S0(dff_q_1)
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(mux_o_370),
  .I1(mux_o_371),
  .S0(dff_q_1)
);
MUX2 mux_inst_374 (
  .O(dout[24]),
  .I0(mux_o_372),
  .I1(mux_o_373),
  .S0(dff_q_0)
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(sp_inst_16_dout[25]),
  .I1(sp_inst_17_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(sp_inst_18_dout[25]),
  .I1(sp_inst_19_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_377 (
  .O(mux_o_377),
  .I0(sp_inst_20_dout[25]),
  .I1(sp_inst_21_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_378 (
  .O(mux_o_378),
  .I0(sp_inst_22_dout[25]),
  .I1(sp_inst_23_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_379 (
  .O(mux_o_379),
  .I0(sp_inst_24_dout[25]),
  .I1(sp_inst_25_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_380 (
  .O(mux_o_380),
  .I0(sp_inst_26_dout[25]),
  .I1(sp_inst_27_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_381 (
  .O(mux_o_381),
  .I0(sp_inst_28_dout[25]),
  .I1(sp_inst_29_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_382 (
  .O(mux_o_382),
  .I0(sp_inst_30_dout[25]),
  .I1(sp_inst_31_dout[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_383 (
  .O(mux_o_383),
  .I0(mux_o_375),
  .I1(mux_o_376),
  .S0(dff_q_2)
);
MUX2 mux_inst_384 (
  .O(mux_o_384),
  .I0(mux_o_377),
  .I1(mux_o_378),
  .S0(dff_q_2)
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(mux_o_379),
  .I1(mux_o_380),
  .S0(dff_q_2)
);
MUX2 mux_inst_386 (
  .O(mux_o_386),
  .I0(mux_o_381),
  .I1(mux_o_382),
  .S0(dff_q_2)
);
MUX2 mux_inst_387 (
  .O(mux_o_387),
  .I0(mux_o_383),
  .I1(mux_o_384),
  .S0(dff_q_1)
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(mux_o_385),
  .I1(mux_o_386),
  .S0(dff_q_1)
);
MUX2 mux_inst_389 (
  .O(dout[25]),
  .I0(mux_o_387),
  .I1(mux_o_388),
  .S0(dff_q_0)
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(sp_inst_16_dout[26]),
  .I1(sp_inst_17_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(sp_inst_18_dout[26]),
  .I1(sp_inst_19_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(sp_inst_20_dout[26]),
  .I1(sp_inst_21_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(sp_inst_22_dout[26]),
  .I1(sp_inst_23_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(sp_inst_24_dout[26]),
  .I1(sp_inst_25_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(sp_inst_26_dout[26]),
  .I1(sp_inst_27_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(sp_inst_28_dout[26]),
  .I1(sp_inst_29_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(sp_inst_30_dout[26]),
  .I1(sp_inst_31_dout[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(mux_o_390),
  .I1(mux_o_391),
  .S0(dff_q_2)
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(mux_o_392),
  .I1(mux_o_393),
  .S0(dff_q_2)
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(mux_o_394),
  .I1(mux_o_395),
  .S0(dff_q_2)
);
MUX2 mux_inst_401 (
  .O(mux_o_401),
  .I0(mux_o_396),
  .I1(mux_o_397),
  .S0(dff_q_2)
);
MUX2 mux_inst_402 (
  .O(mux_o_402),
  .I0(mux_o_398),
  .I1(mux_o_399),
  .S0(dff_q_1)
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(mux_o_400),
  .I1(mux_o_401),
  .S0(dff_q_1)
);
MUX2 mux_inst_404 (
  .O(dout[26]),
  .I0(mux_o_402),
  .I1(mux_o_403),
  .S0(dff_q_0)
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(sp_inst_16_dout[27]),
  .I1(sp_inst_17_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(sp_inst_18_dout[27]),
  .I1(sp_inst_19_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(sp_inst_20_dout[27]),
  .I1(sp_inst_21_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_408 (
  .O(mux_o_408),
  .I0(sp_inst_22_dout[27]),
  .I1(sp_inst_23_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(sp_inst_24_dout[27]),
  .I1(sp_inst_25_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(sp_inst_26_dout[27]),
  .I1(sp_inst_27_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(sp_inst_28_dout[27]),
  .I1(sp_inst_29_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_412 (
  .O(mux_o_412),
  .I0(sp_inst_30_dout[27]),
  .I1(sp_inst_31_dout[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(mux_o_405),
  .I1(mux_o_406),
  .S0(dff_q_2)
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(mux_o_407),
  .I1(mux_o_408),
  .S0(dff_q_2)
);
MUX2 mux_inst_415 (
  .O(mux_o_415),
  .I0(mux_o_409),
  .I1(mux_o_410),
  .S0(dff_q_2)
);
MUX2 mux_inst_416 (
  .O(mux_o_416),
  .I0(mux_o_411),
  .I1(mux_o_412),
  .S0(dff_q_2)
);
MUX2 mux_inst_417 (
  .O(mux_o_417),
  .I0(mux_o_413),
  .I1(mux_o_414),
  .S0(dff_q_1)
);
MUX2 mux_inst_418 (
  .O(mux_o_418),
  .I0(mux_o_415),
  .I1(mux_o_416),
  .S0(dff_q_1)
);
MUX2 mux_inst_419 (
  .O(dout[27]),
  .I0(mux_o_417),
  .I1(mux_o_418),
  .S0(dff_q_0)
);
MUX2 mux_inst_420 (
  .O(mux_o_420),
  .I0(sp_inst_16_dout[28]),
  .I1(sp_inst_17_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_421 (
  .O(mux_o_421),
  .I0(sp_inst_18_dout[28]),
  .I1(sp_inst_19_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(sp_inst_20_dout[28]),
  .I1(sp_inst_21_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(sp_inst_22_dout[28]),
  .I1(sp_inst_23_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(sp_inst_24_dout[28]),
  .I1(sp_inst_25_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(sp_inst_26_dout[28]),
  .I1(sp_inst_27_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_426 (
  .O(mux_o_426),
  .I0(sp_inst_28_dout[28]),
  .I1(sp_inst_29_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(sp_inst_30_dout[28]),
  .I1(sp_inst_31_dout[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(mux_o_420),
  .I1(mux_o_421),
  .S0(dff_q_2)
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(mux_o_422),
  .I1(mux_o_423),
  .S0(dff_q_2)
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(mux_o_424),
  .I1(mux_o_425),
  .S0(dff_q_2)
);
MUX2 mux_inst_431 (
  .O(mux_o_431),
  .I0(mux_o_426),
  .I1(mux_o_427),
  .S0(dff_q_2)
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(mux_o_428),
  .I1(mux_o_429),
  .S0(dff_q_1)
);
MUX2 mux_inst_433 (
  .O(mux_o_433),
  .I0(mux_o_430),
  .I1(mux_o_431),
  .S0(dff_q_1)
);
MUX2 mux_inst_434 (
  .O(dout[28]),
  .I0(mux_o_432),
  .I1(mux_o_433),
  .S0(dff_q_0)
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(sp_inst_16_dout[29]),
  .I1(sp_inst_17_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(sp_inst_18_dout[29]),
  .I1(sp_inst_19_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(sp_inst_20_dout[29]),
  .I1(sp_inst_21_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(sp_inst_22_dout[29]),
  .I1(sp_inst_23_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(sp_inst_24_dout[29]),
  .I1(sp_inst_25_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_440 (
  .O(mux_o_440),
  .I0(sp_inst_26_dout[29]),
  .I1(sp_inst_27_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(sp_inst_28_dout[29]),
  .I1(sp_inst_29_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(sp_inst_30_dout[29]),
  .I1(sp_inst_31_dout[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(mux_o_435),
  .I1(mux_o_436),
  .S0(dff_q_2)
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(mux_o_437),
  .I1(mux_o_438),
  .S0(dff_q_2)
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(mux_o_439),
  .I1(mux_o_440),
  .S0(dff_q_2)
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(mux_o_441),
  .I1(mux_o_442),
  .S0(dff_q_2)
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(mux_o_443),
  .I1(mux_o_444),
  .S0(dff_q_1)
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(mux_o_445),
  .I1(mux_o_446),
  .S0(dff_q_1)
);
MUX2 mux_inst_449 (
  .O(dout[29]),
  .I0(mux_o_447),
  .I1(mux_o_448),
  .S0(dff_q_0)
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(sp_inst_16_dout[30]),
  .I1(sp_inst_17_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(sp_inst_18_dout[30]),
  .I1(sp_inst_19_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(sp_inst_20_dout[30]),
  .I1(sp_inst_21_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_453 (
  .O(mux_o_453),
  .I0(sp_inst_22_dout[30]),
  .I1(sp_inst_23_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(sp_inst_24_dout[30]),
  .I1(sp_inst_25_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(sp_inst_26_dout[30]),
  .I1(sp_inst_27_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(sp_inst_28_dout[30]),
  .I1(sp_inst_29_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(sp_inst_30_dout[30]),
  .I1(sp_inst_31_dout[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(mux_o_450),
  .I1(mux_o_451),
  .S0(dff_q_2)
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(mux_o_452),
  .I1(mux_o_453),
  .S0(dff_q_2)
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(mux_o_454),
  .I1(mux_o_455),
  .S0(dff_q_2)
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(mux_o_456),
  .I1(mux_o_457),
  .S0(dff_q_2)
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(mux_o_458),
  .I1(mux_o_459),
  .S0(dff_q_1)
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(mux_o_460),
  .I1(mux_o_461),
  .S0(dff_q_1)
);
MUX2 mux_inst_464 (
  .O(dout[30]),
  .I0(mux_o_462),
  .I1(mux_o_463),
  .S0(dff_q_0)
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(sp_inst_16_dout[31]),
  .I1(sp_inst_17_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(sp_inst_18_dout[31]),
  .I1(sp_inst_19_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_467 (
  .O(mux_o_467),
  .I0(sp_inst_20_dout[31]),
  .I1(sp_inst_21_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_468 (
  .O(mux_o_468),
  .I0(sp_inst_22_dout[31]),
  .I1(sp_inst_23_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_469 (
  .O(mux_o_469),
  .I0(sp_inst_24_dout[31]),
  .I1(sp_inst_25_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_470 (
  .O(mux_o_470),
  .I0(sp_inst_26_dout[31]),
  .I1(sp_inst_27_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_471 (
  .O(mux_o_471),
  .I0(sp_inst_28_dout[31]),
  .I1(sp_inst_29_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(sp_inst_30_dout[31]),
  .I1(sp_inst_31_dout[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_473 (
  .O(mux_o_473),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(dff_q_2)
);
MUX2 mux_inst_474 (
  .O(mux_o_474),
  .I0(mux_o_467),
  .I1(mux_o_468),
  .S0(dff_q_2)
);
MUX2 mux_inst_475 (
  .O(mux_o_475),
  .I0(mux_o_469),
  .I1(mux_o_470),
  .S0(dff_q_2)
);
MUX2 mux_inst_476 (
  .O(mux_o_476),
  .I0(mux_o_471),
  .I1(mux_o_472),
  .S0(dff_q_2)
);
MUX2 mux_inst_477 (
  .O(mux_o_477),
  .I0(mux_o_473),
  .I1(mux_o_474),
  .S0(dff_q_1)
);
MUX2 mux_inst_478 (
  .O(mux_o_478),
  .I0(mux_o_475),
  .I1(mux_o_476),
  .S0(dff_q_1)
);
MUX2 mux_inst_479 (
  .O(dout[31]),
  .I0(mux_o_477),
  .I1(mux_o_478),
  .S0(dff_q_0)
);
endmodule //Gowin_SP
