//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10 (64-bit)
//Part Number: GW5AST-LV138FPG676AES
//Device: GW5AST-138
//Device Version: B
//Created Time: Thu Jul 25 18:05:25 2024

module Gowin_SP (dout, clk, oce, ce, reset, wre, ad, din, byte_en);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [14:0] ad;
input [31:0] din;
input [3:0] byte_en;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire [15:0] sp_inst_0_dout_w;
wire [15:0] sp_inst_0_dout;
wire [15:0] sp_inst_1_dout_w;
wire [15:0] sp_inst_1_dout;
wire [15:0] sp_inst_2_dout_w;
wire [15:0] sp_inst_2_dout;
wire [15:0] sp_inst_3_dout_w;
wire [15:0] sp_inst_3_dout;
wire [15:0] sp_inst_4_dout_w;
wire [15:0] sp_inst_4_dout;
wire [15:0] sp_inst_5_dout_w;
wire [15:0] sp_inst_5_dout;
wire [15:0] sp_inst_6_dout_w;
wire [15:0] sp_inst_6_dout;
wire [15:0] sp_inst_7_dout_w;
wire [15:0] sp_inst_7_dout;
wire [15:0] sp_inst_8_dout_w;
wire [15:0] sp_inst_8_dout;
wire [15:0] sp_inst_9_dout_w;
wire [15:0] sp_inst_9_dout;
wire [15:0] sp_inst_10_dout_w;
wire [15:0] sp_inst_10_dout;
wire [15:0] sp_inst_11_dout_w;
wire [15:0] sp_inst_11_dout;
wire [15:0] sp_inst_12_dout_w;
wire [15:0] sp_inst_12_dout;
wire [15:0] sp_inst_13_dout_w;
wire [15:0] sp_inst_13_dout;
wire [15:0] sp_inst_14_dout_w;
wire [15:0] sp_inst_14_dout;
wire [15:0] sp_inst_15_dout_w;
wire [15:0] sp_inst_15_dout;
wire [15:0] sp_inst_16_dout_w;
wire [15:0] sp_inst_16_dout;
wire [15:0] sp_inst_17_dout_w;
wire [15:0] sp_inst_17_dout;
wire [15:0] sp_inst_18_dout_w;
wire [15:0] sp_inst_18_dout;
wire [15:0] sp_inst_19_dout_w;
wire [15:0] sp_inst_19_dout;
wire [15:0] sp_inst_20_dout_w;
wire [15:0] sp_inst_20_dout;
wire [15:0] sp_inst_21_dout_w;
wire [15:0] sp_inst_21_dout;
wire [15:0] sp_inst_22_dout_w;
wire [15:0] sp_inst_22_dout;
wire [15:0] sp_inst_23_dout_w;
wire [15:0] sp_inst_23_dout;
wire [15:0] sp_inst_24_dout_w;
wire [15:0] sp_inst_24_dout;
wire [15:0] sp_inst_25_dout_w;
wire [15:0] sp_inst_25_dout;
wire [15:0] sp_inst_26_dout_w;
wire [15:0] sp_inst_26_dout;
wire [15:0] sp_inst_27_dout_w;
wire [15:0] sp_inst_27_dout;
wire [15:0] sp_inst_28_dout_w;
wire [15:0] sp_inst_28_dout;
wire [15:0] sp_inst_29_dout_w;
wire [15:0] sp_inst_29_dout;
wire [15:0] sp_inst_30_dout_w;
wire [15:0] sp_inst_30_dout;
wire [15:0] sp_inst_31_dout_w;
wire [15:0] sp_inst_31_dout;
wire [15:0] sp_inst_32_dout_w;
wire [31:16] sp_inst_32_dout;
wire [15:0] sp_inst_33_dout_w;
wire [31:16] sp_inst_33_dout;
wire [15:0] sp_inst_34_dout_w;
wire [31:16] sp_inst_34_dout;
wire [15:0] sp_inst_35_dout_w;
wire [31:16] sp_inst_35_dout;
wire [15:0] sp_inst_36_dout_w;
wire [31:16] sp_inst_36_dout;
wire [15:0] sp_inst_37_dout_w;
wire [31:16] sp_inst_37_dout;
wire [15:0] sp_inst_38_dout_w;
wire [31:16] sp_inst_38_dout;
wire [15:0] sp_inst_39_dout_w;
wire [31:16] sp_inst_39_dout;
wire [15:0] sp_inst_40_dout_w;
wire [31:16] sp_inst_40_dout;
wire [15:0] sp_inst_41_dout_w;
wire [31:16] sp_inst_41_dout;
wire [15:0] sp_inst_42_dout_w;
wire [31:16] sp_inst_42_dout;
wire [15:0] sp_inst_43_dout_w;
wire [31:16] sp_inst_43_dout;
wire [15:0] sp_inst_44_dout_w;
wire [31:16] sp_inst_44_dout;
wire [15:0] sp_inst_45_dout_w;
wire [31:16] sp_inst_45_dout;
wire [15:0] sp_inst_46_dout_w;
wire [31:16] sp_inst_46_dout;
wire [15:0] sp_inst_47_dout_w;
wire [31:16] sp_inst_47_dout;
wire [15:0] sp_inst_48_dout_w;
wire [31:16] sp_inst_48_dout;
wire [15:0] sp_inst_49_dout_w;
wire [31:16] sp_inst_49_dout;
wire [15:0] sp_inst_50_dout_w;
wire [31:16] sp_inst_50_dout;
wire [15:0] sp_inst_51_dout_w;
wire [31:16] sp_inst_51_dout;
wire [15:0] sp_inst_52_dout_w;
wire [31:16] sp_inst_52_dout;
wire [15:0] sp_inst_53_dout_w;
wire [31:16] sp_inst_53_dout;
wire [15:0] sp_inst_54_dout_w;
wire [31:16] sp_inst_54_dout;
wire [15:0] sp_inst_55_dout_w;
wire [31:16] sp_inst_55_dout;
wire [15:0] sp_inst_56_dout_w;
wire [31:16] sp_inst_56_dout;
wire [15:0] sp_inst_57_dout_w;
wire [31:16] sp_inst_57_dout;
wire [15:0] sp_inst_58_dout_w;
wire [31:16] sp_inst_58_dout;
wire [15:0] sp_inst_59_dout_w;
wire [31:16] sp_inst_59_dout;
wire [15:0] sp_inst_60_dout_w;
wire [31:16] sp_inst_60_dout;
wire [15:0] sp_inst_61_dout_w;
wire [31:16] sp_inst_61_dout;
wire [15:0] sp_inst_62_dout_w;
wire [31:16] sp_inst_62_dout;
wire [15:0] sp_inst_63_dout_w;
wire [31:16] sp_inst_63_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_91;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_104;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_124;
wire mux_o_125;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_164;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_179;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_209;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_224;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_245;
wire mux_o_246;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_251;
wire mux_o_252;
wire mux_o_253;
wire mux_o_254;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_258;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_265;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_269;
wire mux_o_270;
wire mux_o_271;
wire mux_o_272;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_279;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_284;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_299;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_308;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_314;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_321;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_329;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_335;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_349;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_356;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_360;
wire mux_o_361;
wire mux_o_362;
wire mux_o_363;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_370;
wire mux_o_372;
wire mux_o_373;
wire mux_o_374;
wire mux_o_375;
wire mux_o_376;
wire mux_o_377;
wire mux_o_378;
wire mux_o_379;
wire mux_o_380;
wire mux_o_381;
wire mux_o_382;
wire mux_o_383;
wire mux_o_384;
wire mux_o_385;
wire mux_o_386;
wire mux_o_387;
wire mux_o_388;
wire mux_o_389;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_401;
wire mux_o_403;
wire mux_o_404;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_408;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_412;
wire mux_o_413;
wire mux_o_414;
wire mux_o_415;
wire mux_o_416;
wire mux_o_417;
wire mux_o_418;
wire mux_o_419;
wire mux_o_420;
wire mux_o_421;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_426;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_431;
wire mux_o_432;
wire mux_o_434;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_440;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_449;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_453;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_460;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_465;
wire mux_o_466;
wire mux_o_467;
wire mux_o_468;
wire mux_o_469;
wire mux_o_470;
wire mux_o_471;
wire mux_o_472;
wire mux_o_473;
wire mux_o_474;
wire mux_o_475;
wire mux_o_476;
wire mux_o_477;
wire mux_o_478;
wire mux_o_479;
wire mux_o_480;
wire mux_o_481;
wire mux_o_482;
wire mux_o_483;
wire mux_o_484;
wire mux_o_485;
wire mux_o_486;
wire mux_o_487;
wire mux_o_488;
wire mux_o_489;
wire mux_o_490;
wire mux_o_491;
wire mux_o_492;
wire mux_o_493;
wire mux_o_494;
wire mux_o_496;
wire mux_o_497;
wire mux_o_498;
wire mux_o_499;
wire mux_o_500;
wire mux_o_501;
wire mux_o_502;
wire mux_o_503;
wire mux_o_504;
wire mux_o_505;
wire mux_o_506;
wire mux_o_507;
wire mux_o_508;
wire mux_o_509;
wire mux_o_510;
wire mux_o_511;
wire mux_o_512;
wire mux_o_513;
wire mux_o_514;
wire mux_o_515;
wire mux_o_516;
wire mux_o_517;
wire mux_o_518;
wire mux_o_519;
wire mux_o_520;
wire mux_o_521;
wire mux_o_522;
wire mux_o_523;
wire mux_o_524;
wire mux_o_525;
wire mux_o_527;
wire mux_o_528;
wire mux_o_529;
wire mux_o_530;
wire mux_o_531;
wire mux_o_532;
wire mux_o_533;
wire mux_o_534;
wire mux_o_535;
wire mux_o_536;
wire mux_o_537;
wire mux_o_538;
wire mux_o_539;
wire mux_o_540;
wire mux_o_541;
wire mux_o_542;
wire mux_o_543;
wire mux_o_544;
wire mux_o_545;
wire mux_o_546;
wire mux_o_547;
wire mux_o_548;
wire mux_o_549;
wire mux_o_550;
wire mux_o_551;
wire mux_o_552;
wire mux_o_553;
wire mux_o_554;
wire mux_o_555;
wire mux_o_556;
wire mux_o_558;
wire mux_o_559;
wire mux_o_560;
wire mux_o_561;
wire mux_o_562;
wire mux_o_563;
wire mux_o_564;
wire mux_o_565;
wire mux_o_566;
wire mux_o_567;
wire mux_o_568;
wire mux_o_569;
wire mux_o_570;
wire mux_o_571;
wire mux_o_572;
wire mux_o_573;
wire mux_o_574;
wire mux_o_575;
wire mux_o_576;
wire mux_o_577;
wire mux_o_578;
wire mux_o_579;
wire mux_o_580;
wire mux_o_581;
wire mux_o_582;
wire mux_o_583;
wire mux_o_584;
wire mux_o_585;
wire mux_o_586;
wire mux_o_587;
wire mux_o_589;
wire mux_o_590;
wire mux_o_591;
wire mux_o_592;
wire mux_o_593;
wire mux_o_594;
wire mux_o_595;
wire mux_o_596;
wire mux_o_597;
wire mux_o_598;
wire mux_o_599;
wire mux_o_600;
wire mux_o_601;
wire mux_o_602;
wire mux_o_603;
wire mux_o_604;
wire mux_o_605;
wire mux_o_606;
wire mux_o_607;
wire mux_o_608;
wire mux_o_609;
wire mux_o_610;
wire mux_o_611;
wire mux_o_612;
wire mux_o_613;
wire mux_o_614;
wire mux_o_615;
wire mux_o_616;
wire mux_o_617;
wire mux_o_618;
wire mux_o_620;
wire mux_o_621;
wire mux_o_622;
wire mux_o_623;
wire mux_o_624;
wire mux_o_625;
wire mux_o_626;
wire mux_o_627;
wire mux_o_628;
wire mux_o_629;
wire mux_o_630;
wire mux_o_631;
wire mux_o_632;
wire mux_o_633;
wire mux_o_634;
wire mux_o_635;
wire mux_o_636;
wire mux_o_637;
wire mux_o_638;
wire mux_o_639;
wire mux_o_640;
wire mux_o_641;
wire mux_o_642;
wire mux_o_643;
wire mux_o_644;
wire mux_o_645;
wire mux_o_646;
wire mux_o_647;
wire mux_o_648;
wire mux_o_649;
wire mux_o_651;
wire mux_o_652;
wire mux_o_653;
wire mux_o_654;
wire mux_o_655;
wire mux_o_656;
wire mux_o_657;
wire mux_o_658;
wire mux_o_659;
wire mux_o_660;
wire mux_o_661;
wire mux_o_662;
wire mux_o_663;
wire mux_o_664;
wire mux_o_665;
wire mux_o_666;
wire mux_o_667;
wire mux_o_668;
wire mux_o_669;
wire mux_o_670;
wire mux_o_671;
wire mux_o_672;
wire mux_o_673;
wire mux_o_674;
wire mux_o_675;
wire mux_o_676;
wire mux_o_677;
wire mux_o_678;
wire mux_o_679;
wire mux_o_680;
wire mux_o_682;
wire mux_o_683;
wire mux_o_684;
wire mux_o_685;
wire mux_o_686;
wire mux_o_687;
wire mux_o_688;
wire mux_o_689;
wire mux_o_690;
wire mux_o_691;
wire mux_o_692;
wire mux_o_693;
wire mux_o_694;
wire mux_o_695;
wire mux_o_696;
wire mux_o_697;
wire mux_o_698;
wire mux_o_699;
wire mux_o_700;
wire mux_o_701;
wire mux_o_702;
wire mux_o_703;
wire mux_o_704;
wire mux_o_705;
wire mux_o_706;
wire mux_o_707;
wire mux_o_708;
wire mux_o_709;
wire mux_o_710;
wire mux_o_711;
wire mux_o_713;
wire mux_o_714;
wire mux_o_715;
wire mux_o_716;
wire mux_o_717;
wire mux_o_718;
wire mux_o_719;
wire mux_o_720;
wire mux_o_721;
wire mux_o_722;
wire mux_o_723;
wire mux_o_724;
wire mux_o_725;
wire mux_o_726;
wire mux_o_727;
wire mux_o_728;
wire mux_o_729;
wire mux_o_730;
wire mux_o_731;
wire mux_o_732;
wire mux_o_733;
wire mux_o_734;
wire mux_o_735;
wire mux_o_736;
wire mux_o_737;
wire mux_o_738;
wire mux_o_739;
wire mux_o_740;
wire mux_o_741;
wire mux_o_742;
wire mux_o_744;
wire mux_o_745;
wire mux_o_746;
wire mux_o_747;
wire mux_o_748;
wire mux_o_749;
wire mux_o_750;
wire mux_o_751;
wire mux_o_752;
wire mux_o_753;
wire mux_o_754;
wire mux_o_755;
wire mux_o_756;
wire mux_o_757;
wire mux_o_758;
wire mux_o_759;
wire mux_o_760;
wire mux_o_761;
wire mux_o_762;
wire mux_o_763;
wire mux_o_764;
wire mux_o_765;
wire mux_o_766;
wire mux_o_767;
wire mux_o_768;
wire mux_o_769;
wire mux_o_770;
wire mux_o_771;
wire mux_o_772;
wire mux_o_773;
wire mux_o_775;
wire mux_o_776;
wire mux_o_777;
wire mux_o_778;
wire mux_o_779;
wire mux_o_780;
wire mux_o_781;
wire mux_o_782;
wire mux_o_783;
wire mux_o_784;
wire mux_o_785;
wire mux_o_786;
wire mux_o_787;
wire mux_o_788;
wire mux_o_789;
wire mux_o_790;
wire mux_o_791;
wire mux_o_792;
wire mux_o_793;
wire mux_o_794;
wire mux_o_795;
wire mux_o_796;
wire mux_o_797;
wire mux_o_798;
wire mux_o_799;
wire mux_o_800;
wire mux_o_801;
wire mux_o_802;
wire mux_o_803;
wire mux_o_804;
wire mux_o_806;
wire mux_o_807;
wire mux_o_808;
wire mux_o_809;
wire mux_o_810;
wire mux_o_811;
wire mux_o_812;
wire mux_o_813;
wire mux_o_814;
wire mux_o_815;
wire mux_o_816;
wire mux_o_817;
wire mux_o_818;
wire mux_o_819;
wire mux_o_820;
wire mux_o_821;
wire mux_o_822;
wire mux_o_823;
wire mux_o_824;
wire mux_o_825;
wire mux_o_826;
wire mux_o_827;
wire mux_o_828;
wire mux_o_829;
wire mux_o_830;
wire mux_o_831;
wire mux_o_832;
wire mux_o_833;
wire mux_o_834;
wire mux_o_835;
wire mux_o_837;
wire mux_o_838;
wire mux_o_839;
wire mux_o_840;
wire mux_o_841;
wire mux_o_842;
wire mux_o_843;
wire mux_o_844;
wire mux_o_845;
wire mux_o_846;
wire mux_o_847;
wire mux_o_848;
wire mux_o_849;
wire mux_o_850;
wire mux_o_851;
wire mux_o_852;
wire mux_o_853;
wire mux_o_854;
wire mux_o_855;
wire mux_o_856;
wire mux_o_857;
wire mux_o_858;
wire mux_o_859;
wire mux_o_860;
wire mux_o_861;
wire mux_o_862;
wire mux_o_863;
wire mux_o_864;
wire mux_o_865;
wire mux_o_866;
wire mux_o_868;
wire mux_o_869;
wire mux_o_870;
wire mux_o_871;
wire mux_o_872;
wire mux_o_873;
wire mux_o_874;
wire mux_o_875;
wire mux_o_876;
wire mux_o_877;
wire mux_o_878;
wire mux_o_879;
wire mux_o_880;
wire mux_o_881;
wire mux_o_882;
wire mux_o_883;
wire mux_o_884;
wire mux_o_885;
wire mux_o_886;
wire mux_o_887;
wire mux_o_888;
wire mux_o_889;
wire mux_o_890;
wire mux_o_891;
wire mux_o_892;
wire mux_o_893;
wire mux_o_894;
wire mux_o_895;
wire mux_o_896;
wire mux_o_897;
wire mux_o_899;
wire mux_o_900;
wire mux_o_901;
wire mux_o_902;
wire mux_o_903;
wire mux_o_904;
wire mux_o_905;
wire mux_o_906;
wire mux_o_907;
wire mux_o_908;
wire mux_o_909;
wire mux_o_910;
wire mux_o_911;
wire mux_o_912;
wire mux_o_913;
wire mux_o_914;
wire mux_o_915;
wire mux_o_916;
wire mux_o_917;
wire mux_o_918;
wire mux_o_919;
wire mux_o_920;
wire mux_o_921;
wire mux_o_922;
wire mux_o_923;
wire mux_o_924;
wire mux_o_925;
wire mux_o_926;
wire mux_o_927;
wire mux_o_928;
wire mux_o_930;
wire mux_o_931;
wire mux_o_932;
wire mux_o_933;
wire mux_o_934;
wire mux_o_935;
wire mux_o_936;
wire mux_o_937;
wire mux_o_938;
wire mux_o_939;
wire mux_o_940;
wire mux_o_941;
wire mux_o_942;
wire mux_o_943;
wire mux_o_944;
wire mux_o_945;
wire mux_o_946;
wire mux_o_947;
wire mux_o_948;
wire mux_o_949;
wire mux_o_950;
wire mux_o_951;
wire mux_o_952;
wire mux_o_953;
wire mux_o_954;
wire mux_o_955;
wire mux_o_956;
wire mux_o_957;
wire mux_o_958;
wire mux_o_959;
wire mux_o_961;
wire mux_o_962;
wire mux_o_963;
wire mux_o_964;
wire mux_o_965;
wire mux_o_966;
wire mux_o_967;
wire mux_o_968;
wire mux_o_969;
wire mux_o_970;
wire mux_o_971;
wire mux_o_972;
wire mux_o_973;
wire mux_o_974;
wire mux_o_975;
wire mux_o_976;
wire mux_o_977;
wire mux_o_978;
wire mux_o_979;
wire mux_o_980;
wire mux_o_981;
wire mux_o_982;
wire mux_o_983;
wire mux_o_984;
wire mux_o_985;
wire mux_o_986;
wire mux_o_987;
wire mux_o_988;
wire mux_o_989;
wire mux_o_990;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT5 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_0.INIT = 32'h00000001;
LUT5 lut_inst_1 (
  .F(lut_f_1),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_1.INIT = 32'h00000002;
LUT5 lut_inst_2 (
  .F(lut_f_2),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_2.INIT = 32'h00000004;
LUT5 lut_inst_3 (
  .F(lut_f_3),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_3.INIT = 32'h00000008;
LUT5 lut_inst_4 (
  .F(lut_f_4),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_4.INIT = 32'h00000010;
LUT5 lut_inst_5 (
  .F(lut_f_5),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_5.INIT = 32'h00000020;
LUT5 lut_inst_6 (
  .F(lut_f_6),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_6.INIT = 32'h00000040;
LUT5 lut_inst_7 (
  .F(lut_f_7),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_7.INIT = 32'h00000080;
LUT5 lut_inst_8 (
  .F(lut_f_8),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_8.INIT = 32'h00000100;
LUT5 lut_inst_9 (
  .F(lut_f_9),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_9.INIT = 32'h00000200;
LUT5 lut_inst_10 (
  .F(lut_f_10),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_10.INIT = 32'h00000400;
LUT5 lut_inst_11 (
  .F(lut_f_11),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_11.INIT = 32'h00000800;
LUT5 lut_inst_12 (
  .F(lut_f_12),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_12.INIT = 32'h00001000;
LUT5 lut_inst_13 (
  .F(lut_f_13),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_13.INIT = 32'h00002000;
LUT5 lut_inst_14 (
  .F(lut_f_14),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_14.INIT = 32'h00004000;
LUT5 lut_inst_15 (
  .F(lut_f_15),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_15.INIT = 32'h00008000;
LUT5 lut_inst_16 (
  .F(lut_f_16),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_16.INIT = 32'h00010000;
LUT5 lut_inst_17 (
  .F(lut_f_17),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_17.INIT = 32'h00020000;
LUT5 lut_inst_18 (
  .F(lut_f_18),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_18.INIT = 32'h00040000;
LUT5 lut_inst_19 (
  .F(lut_f_19),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_19.INIT = 32'h00080000;
LUT5 lut_inst_20 (
  .F(lut_f_20),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_20.INIT = 32'h00100000;
LUT5 lut_inst_21 (
  .F(lut_f_21),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_21.INIT = 32'h00200000;
LUT5 lut_inst_22 (
  .F(lut_f_22),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_22.INIT = 32'h00400000;
LUT5 lut_inst_23 (
  .F(lut_f_23),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_23.INIT = 32'h00800000;
LUT5 lut_inst_24 (
  .F(lut_f_24),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_24.INIT = 32'h01000000;
LUT5 lut_inst_25 (
  .F(lut_f_25),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_25.INIT = 32'h02000000;
LUT5 lut_inst_26 (
  .F(lut_f_26),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_26.INIT = 32'h04000000;
LUT5 lut_inst_27 (
  .F(lut_f_27),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_27.INIT = 32'h08000000;
LUT5 lut_inst_28 (
  .F(lut_f_28),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_28.INIT = 32'h10000000;
LUT5 lut_inst_29 (
  .F(lut_f_29),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_29.INIT = 32'h20000000;
LUT5 lut_inst_30 (
  .F(lut_f_30),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_30.INIT = 32'h40000000;
LUT5 lut_inst_31 (
  .F(lut_f_31),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_31.INIT = 32'h80000000;
SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[15:0],sp_inst_0_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b01;
defparam sp_inst_0.BIT_WIDTH = 16;
defparam sp_inst_0.BLK_SEL = 3'b001;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h000CD1CF358E71EF002F018C002C11AD020F3590020F35F0A1EF018F2000000D;
defparam sp_inst_0.INIT_RAM_01 = 256'hFD8CE3EC118CFD8C002C102C000C302C002CF9AC118C018011AC51AD000D018C;
defparam sp_inst_0.INIT_RAM_02 = 256'h0000000000000000002080000020BC00F06300230180200C402C418CA06C442C;
defparam sp_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[15:0],sp_inst_1_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_1}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b01;
defparam sp_inst_1.BIT_WIDTH = 16;
defparam sp_inst_1.BLK_SEL = 3'b001;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'h92A8A2A7B2A6C2A5D2A472B482B392B2A2B1B2B0C2AFD2AEE2ADF2AC0055C435;
defparam sp_inst_1.INIT_RAM_01 = 256'h2DA0818D2DA0418D2DA0218D2DA0118D65A0F18D140C42A352A162AB72AA82A9;
defparam sp_inst_1.INIT_RAM_02 = 256'h140040001C00B40024009C002C0068003400E4003C00A4002DA0018D2DA0018D;
defparam sp_inst_1.INIT_RAM_03 = 256'hC2A5D2A472B482B392B2A2B1B2B0C2AFD2AEE2ADF2AC0055040054000DA0018D;
defparam sp_inst_1.INIT_RAM_04 = 256'hBECC008C80766076706180633800C41542A352A162AB72AA82A992A8A2A7B2A6;
defparam sp_inst_1.INIT_RAM_05 = 256'h52C662C572C4C076A076B0614063002080636076706100008C00D0040185BECC;
defparam sp_inst_1.INIT_RAM_06 = 256'h52CC5000B2C092CC72CC0C0087FFB40492CC300C72CC1D8072CC258042CC42C7;
defparam sp_inst_1.INIT_RAM_07 = 256'hB2CC92CC000709A035CC92CE52CDC1AC35CDC2CEB2CD5DCC00070980B1AE92CD;
defparam sp_inst_1.INIT_RAM_08 = 256'h1D8DB2CCA2CD7400A2CC31CC358CB5CE31ADB2CEB2CD62CCB19F92CCB2CC058C;
defparam sp_inst_1.INIT_RAM_09 = 256'h1400818CC18C818C82CC198D240C82CD82CC000C0800C18C31ACC2CDFD8CA2CC;
defparam sp_inst_1.INIT_RAM_0A = 256'hC063A076B0610184000C8C0CA2CCA2CCFD8CA2CC97FF0184818C5D8C818C82CC;
defparam sp_inst_1.INIT_RAM_0B = 256'h72CC33FF0184BECC3FFF34040DAC280CBECD300072C4C076A076B06140630020;
defparam sp_inst_1.INIT_RAM_0C = 256'hE076F06180630020C063A076B0610184000CC59FBECCBECC018C72CC72CC058C;
defparam sp_inst_1.INIT_RAM_0D = 256'h3000B2C0A2CC72CC72CC918C82CC72CB62CA52C942C832C722C612C532C40076;
defparam sp_inst_1.INIT_RAM_0E = 256'h6D8C018C31AC32CD058CB2CC92CC040CE5AC940C8ECD8ECC018C31AC32CDB2CC;
defparam sp_inst_1.INIT_RAM_0F = 256'hB2CCA2CC118CA2CCDBFF0184018CA2CC0180018C31AC918C014C898DADAC4C0D;
defparam sp_inst_1.INIT_RAM_10 = 256'hA2CC6800B2CC058CB2CCA2CC118CA2CC0FFF0184818C018CA2CC9800B2CC058C;
defparam sp_inst_1.INIT_RAM_11 = 256'h0407018CA2CC3000B2CC058CB2CCA2CC118CA2CC13FF018492C528060007018C;
defparam sp_inst_1.INIT_RAM_12 = 256'h92C520060007018CA2CCF800B2CC058CB2CCA2CC118CA2CCDBFF018492C52806;
defparam sp_inst_1.INIT_RAM_13 = 256'h6BFF018492C508060007018CA2CCC000B2CC058CB2CCA2CC118CA2CCA3FF0184;
defparam sp_inst_1.INIT_RAM_14 = 256'h118CA2CC33FF018492C540060007018CA2CC8800B2CC058CB2CCA2CC118CA2CC;
defparam sp_inst_1.INIT_RAM_15 = 256'h3C0092C0B2CC058CB2CC3800B2CC058CB2CCD3FF94045000B2CC058CB2CCA2CC;
defparam sp_inst_1.INIT_RAM_16 = 256'h058CB2CCB2CC058CB2CC92CC31AC418C018C31CC32CE058CB2CC31AD280C92CD;
defparam sp_inst_1.INIT_RAM_17 = 256'h92CD3C0092C0BBFF958DE40C018D31AC32CD058CB2CCD98DC00C018D31AC32CD;
defparam sp_inst_1.INIT_RAM_18 = 256'h32CD058CB2CCB2CC058CB2CC92CC31AC418C018C31CC32CE058CB2CC31AD280C;
defparam sp_inst_1.INIT_RAM_19 = 256'h24000000B7FF94043FFF958DE40C018D31AC32CD058CB2CC5D8DC00C018D31AC;
defparam sp_inst_1.INIT_RAM_1A = 256'hC59F018C31AC32CDB2CCB2CC058CB2CC8FFF01848ECC9BFF34040DAC280C8ECD;
defparam sp_inst_1.INIT_RAM_1B = 256'h818C158CB2CC0000AECC00ACB2C480767076806300208063E076F0610184000C;
defparam sp_inst_1.INIT_RAM_1C = 256'h406330760000042040763076C0630020806370760000018DAECDB2CCF19F818C;
defparam sp_inst_1.INIT_RAM_1D = 256'h2180C18CD80C40763076C0630020406330760000102C040C40763076C0630020;
defparam sp_inst_1.INIT_RAM_1E = 256'h30760000218D040DC18CD80C118D01AD006DC18CD80C018D01AD138DC18CD80C;
defparam sp_inst_1.INIT_RAM_1F = 256'h31AD018C006C0007098031CD240C31AE000CB2CDB2C480767076806300204063;
defparam sp_inst_1.INIT_RAM_20 = 256'h81AD0DADBECDCE0CBECC008C8076707680630020806370760000118DC18CD80C;
defparam sp_inst_1.INIT_RAM_21 = 256'h807660767061806300208063707600000D8D81AD0DADCE0C818D898CBECC018D;
defparam sp_inst_1.INIT_RAM_22 = 256'h818C058CCE0C0000018D81AD41ADCE0C818D018CCE0C8FFF0184BECCBECC008C;
defparam sp_inst_1.INIT_RAM_23 = 256'h40763076C06300208063607670610000F19F058C818C058CCE0C0000F19F118C;
defparam sp_inst_1.INIT_RAM_24 = 256'h0000158D81ADB5CD7C0DCE0C818E158CCE0C158D81AD09ADCE0C818D158CCE0C;
defparam sp_inst_1.INIT_RAM_25 = 256'h818D158CCE0C158D81AD09ADCE0C818D158CCE0C40763076C063002040633076;
defparam sp_inst_1.INIT_RAM_26 = 256'hB2CC72CC52C662C572C4C076B07640630020406330760000158D81AD81ADCE0C;
defparam sp_inst_1.INIT_RAM_27 = 256'h0020C063B076018472CCDD9F52CDFD8D52CC018D81AD62CDB2CD058DB2CC1C00;
defparam sp_inst_1.INIT_RAM_28 = 256'hB2CC040E018DD60C318062CCB2CC72CC698D7C0C72CD62C572C4C076B0764063;
defparam sp_inst_1.INIT_RAM_29 = 256'h018D39ADD60C018E31CCB2CC040E018DD60C9000018DB9ADD60C018E300C31CC;
defparam sp_inst_1.INIT_RAM_2A = 256'h418DB9ADD60C018E300C31CCB2CC040E418DD60C318062CCB2CC818C72CC6800;
defparam sp_inst_1.INIT_RAM_2B = 256'hB07640630020C063B0760000418D39ADD60C018E31CCB2CC040E418DD60C2800;
defparam sp_inst_1.INIT_RAM_2C = 256'h300C31CCB2CC040E118DD60C318062CCB2CC72CC698D7C0C72CD62C572C4C076;
defparam sp_inst_1.INIT_RAM_2D = 256'h72CC6800118D39ADD60C018E31CCB2CC040E118DD60C9000118DB9ADD60C018E;
defparam sp_inst_1.INIT_RAM_2E = 256'hD60C2800518DB9ADD60C018E300C31CCB2CC040E518DD60C318062CCB2CC818C;
defparam sp_inst_1.INIT_RAM_2F = 256'h72C4C076B07640630020C063B0760000518D39ADD60C018E31CCB2CC040E518D;
defparam sp_inst_1.INIT_RAM_30 = 256'h040C0D8D35CDB2CD040EB58C35CDB2CD040E218CD60CB2CC72CC458D7C0C72CD;
defparam sp_inst_1.INIT_RAM_31 = 256'h0D8D35CDB2CD040EB58C35CDB2CD040E618CD60CB2CC818C72CC4400000C4C00;
defparam sp_inst_1.INIT_RAM_32 = 256'h040D818CFFECBECC008C80766076706180630020C063B0760184000C0800040C;
defparam sp_inst_1.INIT_RAM_33 = 256'hA2C5B2C480767076806300208063607670610000AC002084FFC40185BECC018D;
defparam sp_inst_1.INIT_RAM_34 = 256'hB2CC0000B2C48076707680630020806370760000318DB2CC31ADA2CC318DB2CC;
defparam sp_inst_1.INIT_RAM_35 = 256'hB2CC018D81AD030DB2CCB2C48076707680630020806370760000F59FB2CDFD8D;
defparam sp_inst_1.INIT_RAM_36 = 256'h018CD08CB2C072C4C076B07640630020806370760000198D080DB2CC118D800D;
defparam sp_inst_1.INIT_RAM_37 = 256'hA18DB2CC018D81ADB2CDD20CB2CCFD8C898CB2CCB2CCA00C098D800DD20CA2CC;
defparam sp_inst_1.INIT_RAM_38 = 256'h0020C063B0760000118D100DD20C1180198C72CC098D880DD20C058D81ADD20C;
defparam sp_inst_1.INIT_RAM_39 = 256'h806370760000118DFC0DD20C1000118D000DD20C1580B2CCB2C4807670768063;
defparam sp_inst_1.INIT_RAM_3A = 256'h70760000118DFC0DD20C1000118D000DD20C1580B2CCB2C48076707680630020;
defparam sp_inst_1.INIT_RAM_3B = 256'h0000118D400DD20C0D8DBECDD20C7800BECC008C807660767061806300208063;
defparam sp_inst_1.INIT_RAM_3C = 256'hBECCBECC118CD20C1000A2C0BECC118CD20C8076707680630020806360767061;
defparam sp_inst_1.INIT_RAM_3D = 256'hD20C1180118CBECCBECC118CD20C8076707680630020806370760000ED9F098C;
defparam sp_inst_1.INIT_RAM_3E = 256'h406330760000D18DA9ADB4ADD60C40763076C0630020806370760000118D100D;
defparam sp_inst_1.INIT_RAM_3F = 256'h4C0404050FFF480404051BFF3404040527FF0404040580766076706180630020;

SP sp_inst_2 (
    .DO({sp_inst_2_dout_w[15:0],sp_inst_2_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_2}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_2.READ_MODE = 1'b0;
defparam sp_inst_2.WRITE_MODE = 2'b01;
defparam sp_inst_2.BIT_WIDTH = 16;
defparam sp_inst_2.BLK_SEL = 3'b001;
defparam sp_inst_2.RESET_MODE = "SYNC";
defparam sp_inst_2.INIT_RAM_00 = 256'hC7FF94040405D3FF90040405DFFF8C040405EBFF88040405F7FF5004040503FF;
defparam sp_inst_2.INIT_RAM_01 = 256'h00058BFF4004000597FF3C040005A3FF38040005AFFF9C040405BBFF98040005;
defparam sp_inst_2.INIT_RAM_02 = 256'h00000000000000000000000000000000000000008400B2CCC98C0E2C7FFF4404;
defparam sp_inst_2.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_04 = 256'hBFFF94040405CBFF90040405759FB2CDFD8DB2CC000000000000000000000000;
defparam sp_inst_2.INIT_RAM_05 = 256'h000083FF8C0400058FFF9C0404059BFF98040405A7FF34040405B3FF04040405;
defparam sp_inst_2.INIT_RAM_06 = 256'h958C016CF3FF018492CCB7FF018492CC80766076706180630020806360767061;
defparam sp_inst_2.INIT_RAM_07 = 256'h000000000000000000000000000000000000000000000000000000008400B2CC;
defparam sp_inst_2.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_09 = 256'hEFFF807660767061806300208063607670610000759FB2CDFD8DB2CC00000000;
defparam sp_inst_2.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000008400B2CC958C016C;
defparam sp_inst_2.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_0C = 256'h20763061C06300208063607670610000759FB2CDFD8DB2CC0000000000000000;
defparam sp_inst_2.INIT_RAM_0D = 256'h600050008800E800407620763061C063002040632076306100002BFF08044076;
defparam sp_inst_2.INIT_RAM_0E = 256'h2076306100004BFF04040005407620763061C06300204063207630610000A400;
defparam sp_inst_2.INIT_RAM_0F = 256'h70618063002040632076306100001BFF04040405407620763061C06300204063;
defparam sp_inst_2.INIT_RAM_10 = 256'h00000000000000000000000000008400B2CC958C016CEBFF8C04040580766076;
defparam sp_inst_2.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_12 = 256'h3FFF8C040005759FB2CDFD8DB2CC000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000008400A2CC958C016C;
defparam sp_inst_2.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_15 = 256'h0000840092CC958C016C93FF8C040405759FA2CDFD8DA2CC0000000000000000;
defparam sp_inst_2.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_17 = 256'h92CC000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_18 = 256'h0405807660767061806300208063607670610000E7FF8C040005759F92CDFD8D;
defparam sp_inst_2.INIT_RAM_19 = 256'h00000000000000000000000000000000000000008400B2CC798C088CB7FF8C04;
defparam sp_inst_2.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_1B = 256'h6076706100000BFF8C040005759FB2CDFD8DB2CC000000000000000000000000;
defparam sp_inst_2.INIT_RAM_1C = 256'h0405C3FF4C040405CFFF50040405DBFF88040405407620763061C06300208063;
defparam sp_inst_2.INIT_RAM_1D = 256'h8400B2CCD98C008C9FFF807660767061806300204063207630610000B7FF4804;
defparam sp_inst_2.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_20 = 256'h00008400A2CCD98C008C6180008CD3FF3804E3FF48040005759FB2CDFD8DB2CC;
defparam sp_inst_2.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_22 = 256'hA2CC000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_23 = 256'h0000000000000000840092CCD98C008CF59F008C1FFF38040000759FA2CDFD8D;
defparam sp_inst_2.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_25 = 256'h759F92CDFD8D92CC000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_26 = 256'h000000000000000000000000840082CCD98C008C6180008C67FF3C048C00040C;
defparam sp_inst_2.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_28 = 256'h3C040000759F82CDFD8D82CC0000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_29 = 256'h000000000000000000000000000000000000840072CCD98C008CF59F008CB3FF;
defparam sp_inst_2.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_2B = 256'h008CFBFF40042000140C759F72CDFD8D72CC0000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_2C = 256'h00000000000000000000000000000000000000000000840062CCD98C008C6180;
defparam sp_inst_2.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_2E = 256'hD98C008CF59F008C47FF40040000759F62CDFD8D62CC00000000000000000000;
defparam sp_inst_2.INIT_RAM_2F = 256'h00000000000000000000000000000000000000000000000000000000840052CC;
defparam sp_inst_2.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_31 = 256'h840042CCD98C008C6180008C8FFF4404B400240C759F52CDFD8D52CC00000000;
defparam sp_inst_2.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_34 = 256'h000000000000840032CCD98C008CF59F008CDBFF44040000759F42CDFD8D42CC;
defparam sp_inst_2.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_36 = 256'h32CDFD8D32CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_37 = 256'h0000840022CCD98C008C6180008C13FF380423FF4C0400053FFF4800340C759F;
defparam sp_inst_2.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_39 = 256'h22CC000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3A = 256'h0000000000000000840012CCD98C008CF59F008C5FFF38040000759F22CDFD8D;
defparam sp_inst_2.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3C = 256'h759F12CDFD8D12CC000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3D = 256'h000000000000000000000000840002CCD98C008C6180008CA7FF3C04CC00080C;
defparam sp_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3F = 256'h3C040000759F02CDFD8D02CC0000000000000000000000000000000000000000;

SP sp_inst_3 (
    .DO({sp_inst_3_dout_w[15:0],sp_inst_3_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_3}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_3.READ_MODE = 1'b0;
defparam sp_inst_3.WRITE_MODE = 2'b01;
defparam sp_inst_3.BIT_WIDTH = 16;
defparam sp_inst_3.BLK_SEL = 3'b001;
defparam sp_inst_3.RESET_MODE = "SYNC";
defparam sp_inst_3.INIT_RAM_00 = 256'h0000000000000000000000000000000000008400F2CCD98C008CF59F008CF3FF;
defparam sp_inst_3.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_02 = 256'h008C3BFF40046000180C759FF2CDFD8DF2CC0000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_03 = 256'h000000000000000000000000000000000000000000008400E2CCD98C008C6180;
defparam sp_inst_3.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_05 = 256'hD98C008CF59F008C87FF40040000759FE2CDFD8DE2CC00000000000000000000;
defparam sp_inst_3.INIT_RAM_06 = 256'h000000000000000000000000000000000000000000000000000000008400D2CC;
defparam sp_inst_3.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_08 = 256'h8400C2CCD98C008C6180008CCFFF4404F400280C759FD2CDFD8DD2CC00000000;
defparam sp_inst_3.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0B = 256'h0000000000008400B2CCD98C008CF59F008C1BFF44040000759FC2CDFD8DC2CC;
defparam sp_inst_3.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0D = 256'hB2CDFD8DB2CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0E = 256'h00008400A2CCD98C008C6180008C53FF380463FF500400057FFF8800380C759F;
defparam sp_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_10 = 256'hA2CC000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_11 = 256'h0000000000000000840092CCD98C008CF59F008C9FFF38040000759FA2CDFD8D;
defparam sp_inst_3.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_13 = 256'h759F92CDFD8D92CC000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_14 = 256'h000000000000000000000000840082CCD98C008C6180008CE7FF3C040C000C0C;
defparam sp_inst_3.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_16 = 256'h3C040000759F82CDFD8D82CC0000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_17 = 256'h000000000000000000000000000000000000840072CCD98C008CF59F008C33FF;
defparam sp_inst_3.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_19 = 256'h008C7BFF4004A0001C0C759F72CDFD8D72CC0000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1A = 256'h00000000000000000000000000000000000000000000840062CCD98C008C6180;
defparam sp_inst_3.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1C = 256'hD98C008CF59F008CC7FF40040000759F62CDFD8D62CC00000000000000000000;
defparam sp_inst_3.INIT_RAM_1D = 256'h00000000000000000000000000000000000000000000000000000000840052CC;
defparam sp_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1F = 256'h840042CCD98C008C6180008C0FFF440434002C0C759F52CDFD8D52CC00000000;
defparam sp_inst_3.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_22 = 256'h000000000000840032CCD98C008CF59F008C5BFF44040000759F42CDFD8D42CC;
defparam sp_inst_3.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_24 = 256'h32CDFD8D32CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_25 = 256'h0000840022CCD98C008C6180008C93FF3804A3FF88040005BFFFC8003C0C759F;
defparam sp_inst_3.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_27 = 256'h22CC000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_28 = 256'h0000000000000000840012CCD98C008CF59F008CDFFF38040000759F22CDFD8D;
defparam sp_inst_3.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2A = 256'h759F12CDFD8D12CC000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2B = 256'h000000000000000000000000840002CCD98C008C6180008C27FF3C044C00100C;
defparam sp_inst_3.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2D = 256'h3C040000759F02CDFD8D02CC0000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2E = 256'h0000000000000000000000000000000000008400F2CCD98C008CF59F008C73FF;
defparam sp_inst_3.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_30 = 256'h008CBBFF4004E000200C759FF2CDFD8DF2CC0000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_31 = 256'h000000000000000000000000000000000000000000008400E2CCD98C008C6180;
defparam sp_inst_3.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_33 = 256'hD98C008CF59F008C07FF40040000759FE2CDFD8DE2CC00000000000000000000;
defparam sp_inst_3.INIT_RAM_34 = 256'h000000000000000000000000000000000000000000000000000000008400D2CC;
defparam sp_inst_3.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_36 = 256'h8400C2CCD98C008C6180008C4FFF44047400300C759FD2CDFD8DD2CC00000000;
defparam sp_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_39 = 256'h0000000000008400B2CCD98C008CF59F008C9BFF44040000759FC2CDFD8DC2CC;
defparam sp_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3B = 256'hB2CDFD8DB2CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3C = 256'h0404BECC008C807660767061806300208063607670610184000C0800400C759F;
defparam sp_inst_3.INIT_RAM_3D = 256'h0000B3FF500417FF0404ABFF67FF0184BECCBBFF77FF0004C7FF83FFE00403FF;
defparam sp_inst_3.INIT_RAM_3E = 256'h00045BFF17FFE00497FF0404BECC008C80766076706180630020806360767061;
defparam sp_inst_3.INIT_RAM_3F = 256'h80630020806360767061000047FF5004ABFF04043FFFFBFF0184BECC4FFF0BFF;

SP sp_inst_4 (
    .DO({sp_inst_4_dout_w[15:0],sp_inst_4_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_4}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_4.READ_MODE = 1'b0;
defparam sp_inst_4.WRITE_MODE = 2'b01;
defparam sp_inst_4.BIT_WIDTH = 16;
defparam sp_inst_4.BLK_SEL = 3'b001;
defparam sp_inst_4.RESET_MODE = "SYNC";
defparam sp_inst_4.INIT_RAM_00 = 256'h0000000000000000000000000000000000008400B2CC418C16CC807660767061;
defparam sp_inst_4.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_02 = 256'h40046FFF800477FFB804759FB2CDFD8DB2CC0000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_03 = 256'h84042FFFFC0437FF04043FFF000447FF40044FFF000457FF20045FFFC00467FF;
defparam sp_inst_4.INIT_RAM_04 = 256'hC004EFFF5404F7FF0004FFFF4C0407FF90040FFFFC0417FFA0041FFF980427FF;
defparam sp_inst_4.INIT_RAM_05 = 256'h5004AFFF3404B7FF8004BFFF6C04C7FF4804CFFF6804D7FF8804DFFF6404E7FF;
defparam sp_inst_4.INIT_RAM_06 = 256'h818CA2CCA2C5B2C48076607670618063002080636076706100009FFFBC04A7FF;
defparam sp_inst_4.INIT_RAM_07 = 256'h398C818CB2CC37FF0184818C418C818C3D8C818C918CB2CC5BFF0184818CC18C;
defparam sp_inst_4.INIT_RAM_08 = 256'h7ECC008CC076A076B06140630020806360767061000017FF0184818C058C818C;
defparam sp_inst_4.INIT_RAM_09 = 256'h01847ECC1C00A2C0BBFF4004C3FF0004CBFF0184818CC18C818CB2CC6400B2C0;
defparam sp_inst_4.INIT_RAM_0A = 256'hA076B0610000998D1C0CB2CDB2CC058CB2CCE18DFC0CA2CDA2CC058CA2CC13FF;
defparam sp_inst_4.INIT_RAM_0B = 256'hA076B0614063002040632076306100004FFF0004407620763061C0630020C063;
defparam sp_inst_4.INIT_RAM_0C = 256'h52CDD800C58D080DB58D040D4ECCA2C0B2C092C04ECC00EC52C662C572C4C076;
defparam sp_inst_4.INIT_RAM_0D = 256'hB2C02BFF72C462C562CC058C62CC72C0158DF80C72CD92CC818C018C31ACA2CC;
defparam sp_inst_4.INIT_RAM_0E = 256'hB2CDB2CC058CB2CCE7FF0184018C31ACB2CC31AD31CC180C92CEF1AD00ED3C00;
defparam sp_inst_4.INIT_RAM_0F = 256'hA2CC52CD1C004D9F018C31ACA2CC52CDA2CC058CA2CC72CC198C72CCC18D140C;
defparam sp_inst_4.INIT_RAM_10 = 256'h3800B2C06FFF72C462C562CC058C62CC72C0158DE00C72CD92CC818C018C31AC;
defparam sp_inst_4.INIT_RAM_11 = 256'hC58D1C0CB2CDB2CC058CB2CC2FFF0184018C31AC61AD00ED31ACB2CC918D92CC;
defparam sp_inst_4.INIT_RAM_12 = 256'h018C31ACE1AD00ED218C31ACB2CC918D92CC3C00B2C013FF72C40185058C62CC;
defparam sp_inst_4.INIT_RAM_13 = 256'hA2CC52CDA2CC058CA2CC72CC218C72CCC18D1C0CB2CDB2CC058CB2CCCFFF0184;
defparam sp_inst_4.INIT_RAM_14 = 256'h00CC62C572C4C076A076B06140630020C063A076B06100000000F19F018C31AC;
defparam sp_inst_4.INIT_RAM_15 = 256'h0184018C31ACA2CCD1ADFFAD3800BEC047FF72C462C5A2CC958C5ECCBEC05ECC;
defparam sp_inst_4.INIT_RAM_16 = 256'hBEC0EBFF72C40185058C62CCC58D3C0CBECDBECC058CBECCA2CC058CA2CC13FF;
defparam sp_inst_4.INIT_RAM_17 = 256'h3C0CBECDBECC058CBECCA2CC058CA2CCB7FF0184018C31ACA2CC61ADFFAD3800;
defparam sp_inst_4.INIT_RAM_18 = 256'h4800B2C042C752C662C572C4C076A076B06140630020C063A076B0610000C58D;
defparam sp_inst_4.INIT_RAM_19 = 256'h058CB2CCB3FF01C462C50186818C31AC818C52CC818DB2CC31AE72CC918DB2CC;
defparam sp_inst_4.INIT_RAM_1A = 256'h52C662C572C40076E076F06100630020C063A076B0610000B5AC42CCB2CDB2CC;
defparam sp_inst_4.INIT_RAM_1B = 256'h92CC62CC92CC058C8D8C42CC140092CC8D8C42CC15801D8C42CCB2C032C842C7;
defparam sp_inst_4.INIT_RAM_1C = 256'hA2CC5BFF0184018C31AC32CDB2CD058DB2CC3000A2CC72CC97FF72C492C56000;
defparam sp_inst_4.INIT_RAM_1D = 256'h00200063E076F06100009DAC42CC92CD92CC058C92CCCDAC52CCA2CDA2CC058C;
defparam sp_inst_4.INIT_RAM_1E = 256'hA2CC818C5ECCB2C0A2C05ACC01AC5ECC00ED00CC62C572C4C076A076B0614063;
defparam sp_inst_4.INIT_RAM_1F = 256'hA2CC3800B2C0B3FF72C462C5BDAC400C5ACD62CC098C62CC72C0158DFC0C72CD;
defparam sp_inst_4.INIT_RAM_20 = 256'h62CCC58D1C0CB2CDB2CC058CB2CC73FF0184018C31AC71AD00ED31ACB2CC918D;
defparam sp_inst_4.INIT_RAM_21 = 256'h0184018C31ACF1AD00ED218C31ACB2CC918DA2CC3C00B2C057FF72C40185058C;
defparam sp_inst_4.INIT_RAM_22 = 256'hA2CE31AD00CD3C00B2C0FBFF72C462C55C00C18D1C0CB2CDB2CC058CB2CC13FF;
defparam sp_inst_4.INIT_RAM_23 = 256'hB0610000C18D140CB2CDB2CC058CB2CCB7FF0184018C31ACB2CC31AD31CC180C;
defparam sp_inst_4.INIT_RAM_24 = 256'h62CCB2CC31AC72CCB2CD1400B2CC040C62C572C4C076B07640630020C063A076;
defparam sp_inst_4.INIT_RAM_25 = 256'h00EC52C662C572C4C076A076B06140630020C063B0760184B2CCE59F62CDFD8D;
defparam sp_inst_4.INIT_RAM_26 = 256'h52CC008D5BFF28040185FD8C31ACB2CC4ECD0400B2C0A2C04ACC01AC4ECC010D;
defparam sp_inst_4.INIT_RAM_27 = 256'h92CC518DB2CC018DFD8C4ECC6580A2CC92CC000709A0B5CC280D000709A0358E;
defparam sp_inst_4.INIT_RAM_28 = 256'h54004BFF018462C5800601A74ACD31AC72CC31ADB2CC018D818C858C4ACC4180;
defparam sp_inst_4.INIT_RAM_29 = 256'h01C74ACE818CC18C818C92CC31AD72CC31ADB2CC018D818C858C4ACCA2CC040C;
defparam sp_inst_4.INIT_RAM_2A = 256'h40630020C063A076B0610000F9ACB2CD4ECCB2CC058CB2CCF7FF01A462C50186;
defparam sp_inst_4.INIT_RAM_2B = 256'h1C0092CC62CCA2CCB2CC8C0072CC8580018C62CCB2CC72CC62C572C4C076B076;
defparam sp_inst_4.INIT_RAM_2C = 256'h018C92CC018DA2CC1980018C92CC2580018CA2CC92CC058C92CCA2CC058CA2CC;
defparam sp_inst_4.INIT_RAM_2D = 256'hC063B0760184000C819F018CB2CCB2CC058CB2CC2000B2CC0D80018C92CCC1AC;
defparam sp_inst_4.INIT_RAM_2E = 256'h0000018DBECDD00CF19F818C818C158CD00C0000BECC008C8076707680630020;
defparam sp_inst_4.INIT_RAM_2F = 256'h8BFF040493FFBC04B7FFA084FF8400054006407620763061C063002080637076;
defparam sp_inst_4.INIT_RAM_30 = 256'h4BFF0184818CE18C018CE18CFFAC407620763061C06300204063207630610000;
defparam sp_inst_4.INIT_RAM_31 = 256'h918CFFAC13FF0184818CA18C018C018CFFAC2FFF0184818CC18C018C718CFFAC;
defparam sp_inst_4.INIT_RAM_32 = 256'hBECCBECC008C807660767061806300204063207630610000FBFF0184818C018C;
defparam sp_inst_4.INIT_RAM_33 = 256'h0184818CA18CB2CCB2C4807660767061806300208063607670610000C3FF0184;
defparam sp_inst_4.INIT_RAM_34 = 256'hBECC008C80766076706180630020806360767061000077FF0184818CB2CC87FF;
defparam sp_inst_4.INIT_RAM_35 = 256'hA18CBACCBACC008C8076607670618063002080636076706100003FFF0184BECC;
defparam sp_inst_4.INIT_RAM_36 = 256'h60767061806300208063607670610000EBFF0184818CBACCFBFF0184818C818C;
defparam sp_inst_4.INIT_RAM_37 = 256'h31ACA2CCC1ADFFAD2C00A2C033FFEFFF258D040DF18CFF8CB2CC418C004C8076;
defparam sp_inst_4.INIT_RAM_38 = 256'h92C0F19F058C818C158CD00C0000D18D240CA2CDA2CC058CA2CC7FFF0184018C;
defparam sp_inst_4.INIT_RAM_39 = 256'hD00C1800098D81AD35CDF40DD00C818E098CD00C2980B2CCB2CCFD8CB2CCA800;
defparam sp_inst_4.INIT_RAM_3A = 256'hFF8E818D018CD00C2400018031AC92CCD1ADFF8D1D80B2CCB99F058C818C158C;
defparam sp_inst_4.INIT_RAM_3B = 256'h258C618CFF8C8D8D2C0C92CD92CC058C92CCB2CCC18C00EC018D31CC92CC41CE;
defparam sp_inst_4.INIT_RAM_3C = 256'h7BFFC4000804407620763061C06300208063607670610184040C0800000C0D80;
defparam sp_inst_4.INIT_RAM_3D = 256'h72CCBC0CB2CC3ACC3ACC008C0076E076F061006300204063207630610184008C;
defparam sp_inst_4.INIT_RAM_3E = 256'h918CFFAC7ECC818CC18C018CF18CFFAC7ACC818CE18C018C518CFFAC76CC040C;
defparam sp_inst_4.INIT_RAM_3F = 256'h818C158CD00C00008EC08ACC1C0C86CC818C018C318CFFAC82CC818CA18C018C;

SP sp_inst_5 (
    .DO({sp_inst_5_dout_w[15:0],sp_inst_5_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_5}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_5.READ_MODE = 1'b0;
defparam sp_inst_5.WRITE_MODE = 2'b01;
defparam sp_inst_5.BIT_WIDTH = 16;
defparam sp_inst_5.BLK_SEL = 3'b001;
defparam sp_inst_5.RESET_MODE = "SYNC";
defparam sp_inst_5.INIT_RAM_00 = 256'h81AD35CDF40DD00C818E098CD00C2980B2CCB2CCFD8CB2CCC000A2C0F19F058C;
defparam sp_inst_5.INIT_RAM_01 = 256'hD00C2400018031ACA2CCA1ADFF8D1D80B2CCB99F058C818C158CD00C1800098D;
defparam sp_inst_5.INIT_RAM_02 = 256'hB2CC3ACC00000184018C31ACA2CCC1ADFF8D018D31CCA2CC11CEFF8E818D018C;
defparam sp_inst_5.INIT_RAM_03 = 256'h080092CC0D8092CC92C4D7FFB084FF84018572CC758D600CA2CDA2CC058CA2CC;
defparam sp_inst_5.INIT_RAM_04 = 256'hA3FF0C0473FF0404EBFFA7FF807660767061806300200063E076F0610184000C;
defparam sp_inst_5.INIT_RAM_05 = 256'hBECC258CA2CC1580A2CCA2C4F7FF4184004C0BFF0184B2CCB2CC140CE7FF0404;
defparam sp_inst_5.INIT_RAM_06 = 256'h13FF7ECC008CC076A076B061406300208063607670610184BECCBECCFC0C0C00;
defparam sp_inst_5.INIT_RAM_07 = 256'h0184B2CCB2CC1D8C818C7ECCA3FF01847ECC53FF08040FFF1004DFFF040457FF;
defparam sp_inst_5.INIT_RAM_08 = 256'hB0610184BECCBECCFC0C0C00BECC258CA2CC1580A2CCA2C44FFF4184004C63FF;
defparam sp_inst_5.INIT_RAM_09 = 256'h1C0CB3FF0C046FFF0C043FFF0404B7FF73FF80766076706180630020C063A076;
defparam sp_inst_5.INIT_RAM_0A = 256'hBECCFC0C0C00BECC258CA2CC1580A2CCA2C4C3FF4184004CD7FF0184B2CCB2CC;
defparam sp_inst_5.INIT_RAM_0B = 256'hE3FF0C04B3FF04042BFFE7FF807660767061806300208063607670610184BECC;
defparam sp_inst_5.INIT_RAM_0C = 256'hBECC258CA2CC1580A2CCA2C437FF4184004C4BFF0184B2CCB2CC240C27FF1404;
defparam sp_inst_5.INIT_RAM_0D = 256'h7ECC00AD008CC076A076B061406300208063607670610184BECCBECCFC0C0C00;
defparam sp_inst_5.INIT_RAM_0E = 256'h818CA18C72CCD7FF01847ECC87FF180443FF180413FF04048BFF47FF72CC01AC;
defparam sp_inst_5.INIT_RAM_0F = 256'h818D31AC818C818C818CA18C72CC818D7ECCAFFF0184818C72CCBFFF0184818C;
defparam sp_inst_5.INIT_RAM_10 = 256'h1580A2CCA2C42BFF4184004C3FFF0184B2CCB2CC358C818C31AC818C818C72CC;
defparam sp_inst_5.INIT_RAM_11 = 256'h80766076706180630020C063A076B0610184BECCBECCFC0C0C00BECC258CA2CC;
defparam sp_inst_5.INIT_RAM_12 = 256'h9FFF4184004CB3FF0184B2CCB2CC440C8FFF34044BFF0C041BFF040493FF4FFF;
defparam sp_inst_5.INIT_RAM_13 = 256'h406300208063607670610184BECCBECCFC0C0C00BECC258CA2CC1580A2CCA2C4;
defparam sp_inst_5.INIT_RAM_14 = 256'h6BFF0404E3FF9FFF6ACC01AC72CC01CC7ECC52C700CD00AE008CC076A076B061;
defparam sp_inst_5.INIT_RAM_15 = 256'h0184818C72CC17FF0184818C818CA18C72CC2FFF01847ECCDFFF6C049BFF2004;
defparam sp_inst_5.INIT_RAM_16 = 256'h818CA18C72CC818D7ECCDFFF0184818C6ACCEFFF0184818C818CA18C6ACC07FF;
defparam sp_inst_5.INIT_RAM_17 = 256'h31AC818C818C6ACC818D31AC818CA18C6ACC818D31AC818C818C72CC818D31AC;
defparam sp_inst_5.INIT_RAM_18 = 256'hA2CCBECC258CA2CC8580A2CCA2C43BFF4184004C4FFF0184B2CCB2CC918C818C;
defparam sp_inst_5.INIT_RAM_19 = 256'h018C318CA2CC018D52CC818D31AC818C018C2D8CA2CC818DA18C818C018C298C;
defparam sp_inst_5.INIT_RAM_1A = 256'h0184BECCBECCFC0C0C00098D52CC818D31AC818C018C358CA2CC818DA18C818C;
defparam sp_inst_5.INIT_RAM_1B = 256'h1FFF78040805F8060807E3FF7ECC008CC076A076B06140630020C063A076B061;
defparam sp_inst_5.INIT_RAM_1C = 256'h00000000000000000000000000008400B2CC918C1C6C0BFFF804080518060807;
defparam sp_inst_5.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_1E = 256'hA076B0610000759FB2CDFD8DB2CC000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_1F = 256'hB6CC49AC140CBACDBACC058CBACCB2C0B6C0BAC0C076A076B06140630020C063;
defparam sp_inst_5.INIT_RAM_20 = 256'hC98C0E2CE7FF78040805E8061007ABFF0180018C31AC718C00CC898D99AC100D;
defparam sp_inst_5.INIT_RAM_21 = 256'h000000000000000000000000000000000000000000000000000000008400A2CC;
defparam sp_inst_5.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_23 = 256'h6ECC6ECC008CB7FF040469806ECC6ECC008C43FF759FA2CDFD8DA2CC00000000;
defparam sp_inst_5.INIT_RAM_24 = 256'h6000B6CC040CBAC0EFFF200408053406040703FFA0040805F8060807C7FF4180;
defparam sp_inst_5.INIT_RAM_25 = 256'h34060407A7FFA0040805F80608076BFF40007BFF01846ECC50008BFF01846ECC;
defparam sp_inst_5.INIT_RAM_26 = 256'h080713FF41806ECC6ECC008C03FF080469806ECC6ECC008C8FFF93FF20040805;
defparam sp_inst_5.INIT_RAM_27 = 256'hD7FF01846ECCAC00B6CC080CBAC03BFF20040805340604074FFFA0040805F806;
defparam sp_inst_5.INIT_RAM_28 = 256'hDFFF2004080534060407F3FFA0040805F8060807B7FF8C00C7FF01846ECC9C00;
defparam sp_inst_5.INIT_RAM_29 = 256'h9FFF2004080534060407B3FFA0040805F806080777FF69806ECC6ECC008C0FFF;
defparam sp_inst_5.INIT_RAM_2A = 256'h080713FFE800B6CC0C0C73FFF80408050806080787FF78040805F80608074BFF;
defparam sp_inst_5.INIT_RAM_2B = 256'hE58C070CA800B6C0E7FF01846ECC3BFFF8040805100608074FFF78040805F806;
defparam sp_inst_5.INIT_RAM_2C = 256'h00000000000000000000000000000000000000000000000000000000840092CC;
defparam sp_inst_5.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_2E = 256'h6ECCB6C0E800B6CC100C11806ECC6ECC008C43FF759F92CDFD8D92CC00000000;
defparam sp_inst_5.INIT_RAM_2F = 256'hB2CC1180B2CCBEC01DAC340CBECDBECC008C87FF9000B2CC040CD4000FFF0184;
defparam sp_inst_5.INIT_RAM_30 = 256'h1005C0C600C60807B2CC058CB2CC118D1C0CB2CDBEC021AC380CBECDB2CCFD8C;
defparam sp_inst_5.INIT_RAM_31 = 256'h0185818CB2CCBEC06DAC3C0CBECD03FFF0041005018604074008B2CCB3FF8004;
defparam sp_inst_5.INIT_RAM_32 = 256'h1005C0C600C608076FFF28040805F806180733FFF5806ECC6ECC008CE3FF0804;
defparam sp_inst_5.INIT_RAM_33 = 256'h000000000000840082CC598C2AAC83FFF0041005018604074008B2CC33FF8004;
defparam sp_inst_5.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_35 = 256'h82CDFD8D82CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_36 = 256'h00000000000000000000840072CCE58C070C00003FFF01846ECCB6C0C000759F;
defparam sp_inst_5.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_38 = 256'hABFF759F72CDFD8D72CC00000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_39 = 256'h9FFF78040805E806100763FFBEC0C076A076B06140630020C063A076B0610000;
defparam sp_inst_5.INIT_RAM_3A = 256'h7ECC7ECC008CF7FF0404D99F7ECC85AC280CBECDBECC058CBECC7ECC008C9BFF;
defparam sp_inst_5.INIT_RAM_3B = 256'h33FF8C0080002004DFFF6D807ECC7ECC008C27FF040400058C06018762CC4980;
defparam sp_inst_5.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000008400A2CCE58C472C;
defparam sp_inst_5.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_3E = 256'h840092CCE58C472CC80024040C008FFF759FA2CDFD8DA2CC0000000000000000;
defparam sp_inst_5.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_6 (
    .DO({sp_inst_6_dout_w[15:0],sp_inst_6_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_6}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_6.READ_MODE = 1'b0;
defparam sp_inst_6.WRITE_MODE = 2'b01;
defparam sp_inst_6.BIT_WIDTH = 16;
defparam sp_inst_6.BLK_SEL = 3'b001;
defparam sp_inst_6.RESET_MODE = "SYNC";
defparam sp_inst_6.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_01 = 256'h000000000000840082CC918C1C6C9BFF1800180477FFD800759F92CDFD8D92CC;
defparam sp_inst_6.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_03 = 256'h82CDFD8D82CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_04 = 256'h80630020C063A076B0610000000063FFFFFF78040805E8061007C3FF2400759F;
defparam sp_inst_6.INIT_RAM_05 = 256'hB2CC918C1C6C63FF0184AECC10009BFF0D80AECCAECC008C27FF807660767061;
defparam sp_inst_6.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000008400;
defparam sp_inst_6.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_08 = 256'hB2C4B2C4807660767061806300208063607670610000759FB2CDFD8DB2CC0000;
defparam sp_inst_6.INIT_RAM_09 = 256'h4063207630610000BFFF0004407620763061C063002080636076706100008BFF;
defparam sp_inst_6.INIT_RAM_0A = 256'h407620763061C0630020406320763061000093FF5404407620763061C0630020;
defparam sp_inst_6.INIT_RAM_0B = 256'h00008400B2CC958C016C80766076706180630020406320763061000067FF0004;
defparam sp_inst_6.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0D = 256'hB2CC000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0E = 256'h000000000000000000000000000000008400A2CCED8C004CFC00759FB2CDFD8D;
defparam sp_inst_6.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_10 = 256'h92CCED8C004C5800759FA2CDFD8DA2CC00000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000008400;
defparam sp_inst_6.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_13 = 256'h000000000000000000000000840082CCED8C004C2C00759F92CDFD8D92CC0000;
defparam sp_inst_6.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_15 = 256'h00008400759F82CDFD8D82CC0000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_16 = 256'h5D8DF98C5D8C858C7ECCAEC07ECC008CC076A076B06140630020806360767061;
defparam sp_inst_6.INIT_RAM_17 = 256'hCE0C0000F19F118C818C058CCE0C0000098DAACDCE0C27FFAACC5D8C31AC000C;
defparam sp_inst_6.INIT_RAM_18 = 256'h0000F19F118C818C058CCE0C00000980CE0CAECC098CCE0CF19F058C818C058C;
defparam sp_inst_6.INIT_RAM_19 = 256'h00000000000000008400B2CC080CEFFFAECC098CCE0CF19F058C818C058CCE0C;
defparam sp_inst_6.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_1B = 256'h759FB2CDFD8DB2CC000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_1C = 256'h7ECC7ACC01AC7ECC00AD008CC076A076B06140630020C063A076B0610184AECC;
defparam sp_inst_6.INIT_RAM_1D = 256'hCE0C0000F19F118C818C058CCE0C0000098DAECDCE0CA7FFAECCF98C818C858C;
defparam sp_inst_6.INIT_RAM_1E = 256'hF19F118C818C058CCE0C0000098D7ACDCE0CAACC098CCE0CF19F058C818C058C;
defparam sp_inst_6.INIT_RAM_1F = 256'h0000000000008400B2CC080C6BFFAACC098CCE0CF19F058C818C058CCE0C0000;
defparam sp_inst_6.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_21 = 256'hB2CDFD8DB2CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_22 = 256'hBEC07ACC01AC7ECC00AD008CC076A076B06140630020C063A076B0610000759F;
defparam sp_inst_6.INIT_RAM_23 = 256'hB061000027FF018401A57ECC818D5D8C31ACBECC7ACDBECC008CCBFF01847ECC;
defparam sp_inst_6.INIT_RAM_24 = 256'h57FF01847ECCBEC07ACC01AC7ECC00AD008CC076A076B06140630020C063A076;
defparam sp_inst_6.INIT_RAM_25 = 256'hA076B0610000ABFF018401A57ECC818D5D8CB1ACBECC5D8D300C7ACCBECC008C;
defparam sp_inst_6.INIT_RAM_26 = 256'h00000000000000008400B2CC880C5BFF9404040580766076706180630020C063;
defparam sp_inst_6.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_28 = 256'h759FB2CDFD8DB2CC000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_29 = 256'h00000000000000000000000000000000000000008400A2CC880CB3FF94040005;
defparam sp_inst_6.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2B = 256'h1FFF04043C050BFF94040405759FA2CDFD8DA2CC000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000840092CC880C;
defparam sp_inst_6.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2E = 256'h5FFFB00400056BFFB404780577FF4404F405759F92CDFD8D92CC000000000000;
defparam sp_inst_6.INIT_RAM_2F = 256'h806300208063607670610184000C3BFF5404000547FFAC04F80553FFA8043405;
defparam sp_inst_6.INIT_RAM_30 = 256'h00000000000000000000000000008400B2CC980C07FF54040005807660767061;
defparam sp_inst_6.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_32 = 256'h008CDBFF5004759FB2CDFD8DB2CC000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_33 = 256'h00208063607670610000AECC008CB3FF5404C3FF50040C0511800D8CAECCAECC;
defparam sp_inst_6.INIT_RAM_34 = 256'h9077A076B061406300204063207630610000F7FF50040C05407620763061C063;
defparam sp_inst_6.INIT_RAM_35 = 256'h218D300D7ECCB6C0BAC0BECCF80C7ACC01AC7ECC42C852C700CD62C5008CC076;
defparam sp_inst_6.INIT_RAM_36 = 256'h31AC000CBACD00000800B6CCC00CBACCDC0C1C00B6CC400CBACC480C2D8D380D;
defparam sp_inst_6.INIT_RAM_37 = 256'hA2CC2C00A2C0ABFF2804000537FF0404000537FF100400054FFF08040185818C;
defparam sp_inst_6.INIT_RAM_38 = 256'hDFFF040401857ECCD1ACA2CD7ACCA2CC058CA2CC07FF24040185018C31AC62CD;
defparam sp_inst_6.INIT_RAM_39 = 256'hA2CCFD8CA2CCB2CC008C2BFF1004A2CC018C026C47FF3404000511AC300C7ECD;
defparam sp_inst_6.INIT_RAM_3A = 256'h18041180A2CC5FFF34040005C19F818CB1ACB6CCB2CD1980058CB2CC2580A2CC;
defparam sp_inst_6.INIT_RAM_3B = 256'hCDAC300C7ECDBECCFC0C0D80058C818CB1ACBACCB2CDBEC0F5806D8C008CD3FF;
defparam sp_inst_6.INIT_RAM_3C = 256'h31AD9ECC8D8DFD8CB2CC25809ECC9ECC1D8C008C7FFF3004B2CC008C8FFF2804;
defparam sp_inst_6.INIT_RAM_3D = 256'hB2CC480C0D8D480CB2CDB2CC040C0D80B2CC018D42CC8D8DB2CC1400018D42CC;
defparam sp_inst_6.INIT_RAM_3E = 256'h0C00D1ACA2CDB2CCA2CC058CA2CC02EC008CFBFF240431B752CDA2CC2C00A2C0;
defparam sp_inst_6.INIT_RAM_3F = 256'h00630020C0639077A076B0610184BECC3FFF04040005CBFF30040005BECCF80C;

SP sp_inst_7 (
    .DO({sp_inst_7_dout_w[15:0],sp_inst_7_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_7}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_7.READ_MODE = 1'b0;
defparam sp_inst_7.WRITE_MODE = 2'b01;
defparam sp_inst_7.BIT_WIDTH = 16;
defparam sp_inst_7.BLK_SEL = 3'b001;
defparam sp_inst_7.RESET_MODE = "SYNC";
defparam sp_inst_7.INIT_RAM_00 = 256'h3ECC63FF50040C05EFFF34041C05EFFF200420053ECC22C5008C0076E076F061;
defparam sp_inst_7.INIT_RAM_01 = 256'h400CA2CD3180BECCBECC008CCFFF30040185040601A701C852CC52CDA2CE52CC;
defparam sp_inst_7.INIT_RAM_02 = 256'h0063E076F0610184BECCBECCF80C0C00018D56CD058C22CC018D22CC52CD25AC;
defparam sp_inst_7.INIT_RAM_03 = 256'h13FF380400052BFF340400052BFF20042005B6C032C40076E076F06100630020;
defparam sp_inst_7.INIT_RAM_04 = 256'hBECCBECC008C03FF30040185080601A701C852CC52CDA2CE56CC800C52CC4C0C;
defparam sp_inst_7.INIT_RAM_05 = 256'hB6CC918D31ACC2CDBACC018D91AD39ADC2CD31AC32CDBACCBACE4C00BAC08180;
defparam sp_inst_7.INIT_RAM_06 = 256'hBECCF80C0DACB6CD918C31ACC2CDBACCB18D0C0CBACDBACC058CBACCB6CCB1AC;
defparam sp_inst_7.INIT_RAM_07 = 256'h30A5FF45BAC0807660767061806300200063E076F0610184BECCD3FF38040005;
defparam sp_inst_7.INIT_RAM_08 = 256'h280C818D818C918C018CB18CFF4C4980008CAFFF0084FF445D80008CFBFF4804;
defparam sp_inst_7.INIT_RAM_09 = 256'h00208063607670610184BACCBACC31AC818C3D8C818C018C218CFF4C818D31AC;
defparam sp_inst_7.INIT_RAM_0A = 256'h0184B2CCB2C00800B2CC040C1180B1AC72CC018DDA0CB2C072C4C076B0764063;
defparam sp_inst_7.INIT_RAM_0B = 256'h018C0D8CD40C018D35CDB2CDDA0C018EDA0CB2C48076707680630020C063B076;
defparam sp_inst_7.INIT_RAM_0C = 256'hD18CFF4C72C4C076B07640630020806370760000018D81AD05AD0D8CD40C818D;
defparam sp_inst_7.INIT_RAM_0D = 256'hD00C058D81ADD00CA18DB2CC0D8D000DD00CB2CCFD8C000709A035CC72CD018E;
defparam sp_inst_7.INIT_RAM_0E = 256'h8076707680630020C063B07600000D8D0C0DD00C098D180DD00C018D81ADB2CD;
defparam sp_inst_7.INIT_RAM_0F = 256'h80630020806370760000018DBECDD00CF19F818C818C158CD00C0000BECC008C;
defparam sp_inst_7.INIT_RAM_10 = 256'h098D81ADFDADD00C818D098CD00CBECC0C0C0D8D0C0CBECDBECC008C80767076;
defparam sp_inst_7.INIT_RAM_11 = 256'h0020806370760000098D81ADD00C5D8D31AC5D8C998CBECC5D8D818C098CD00C;
defparam sp_inst_7.INIT_RAM_12 = 256'h058D318CB2CC018DAECD358C31ADB2CD018CB2CCAECC00ACB2C4807670768063;
defparam sp_inst_7.INIT_RAM_13 = 256'h418DB2CC418DB2CC058D418CB2CC3180B2CC0DAC118CB2CC318DB2CC318DB2CC;
defparam sp_inst_7.INIT_RAM_14 = 256'h118CB2CC218DB2CC218DB2CC058D218CB2CC418DB2CC118DB2CC458D118CB2CC;
defparam sp_inst_7.INIT_RAM_15 = 256'h01CCBFFF1FFFFFFF5BFF807660767061806300208063707600002180B2CC0DAC;
defparam sp_inst_7.INIT_RAM_16 = 256'h00000000000000000000000000000000000000008400B2CCC98C0E2CA7FF0184;
defparam sp_inst_7.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_18 = 256'h00008400A2CCC98C0E2C3BFF759FB2CDFD8DB2CC000000000000000000000000;
defparam sp_inst_7.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_1A = 256'hA2CC000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_1B = 256'hFF2C018D008C6FFFAFFF0180298CFF2CADAC040C008D23FF9804759FA2CDFD8D;
defparam sp_inst_7.INIT_RAM_1C = 256'h018D918CFF4C0180018C31AC018C008C898DBDAC4C0D018C458CFF4C018DB58C;
defparam sp_inst_7.INIT_RAM_1D = 256'h018D080DA58CFF4C29AC340C018D358CFF2C0180218CFF4C2800040419AC040C;
defparam sp_inst_7.INIT_RAM_1E = 256'h818CFF4C018D200DC58CFF4C39AC380C018D558CFF2C4C00018D080D618CFF4C;
defparam sp_inst_7.INIT_RAM_1F = 256'h018DD58CFF2C0180C18CFF4C9000080419AC080C018D318CFF4C1400018D200D;
defparam sp_inst_7.INIT_RAM_20 = 256'h29AC300C018DF58CFF2CBC00018D0C0D018CFF4C018D0C0D458CFF4C29AC2C0C;
defparam sp_inst_7.INIT_RAM_21 = 256'h858CFF4C29AC3C0C018D158CFF2C8400018D100D218CFF4C018D100D658CFF4C;
defparam sp_inst_7.INIT_RAM_22 = 256'h018D040DA58CFF4C39AC400C018D358CFF2C4C00018D3C0D418CFF4C018D3C0D;
defparam sp_inst_7.INIT_RAM_23 = 256'h6C000180A18CFF4C8800100419AC0C0C018D118CFF4C1400018D040D618CFF4C;
defparam sp_inst_7.INIT_RAM_24 = 256'h818CFF4CB800018D080DD18CFF4C018D080D158CFF4CDDAC400C018DA58CFF2C;
defparam sp_inst_7.INIT_RAM_25 = 256'h858CFF4C81AC400C018D158CFF2CAC000180118CFF4C2400140419AC100C018D;
defparam sp_inst_7.INIT_RAM_26 = 256'h818CFF4CC0000C0419AC140C018DF18CFF4C5C00018D080D418CFF4C018D080D;
defparam sp_inst_7.INIT_RAM_27 = 256'hFF2C0400018D180DC18CFF4C018D180D058CFF4C29AC2C0C018D958CFF2C0180;
defparam sp_inst_7.INIT_RAM_28 = 256'h018DD58CFF2CCC00018D1C0DE18CFF4C018D1C0D258CFF4C29AC300C018DB58C;
defparam sp_inst_7.INIT_RAM_29 = 256'h81AC400C018DF58CFF2C9400018D400D018CFF4C018D400D458CFF4C29AC3C0C;
defparam sp_inst_7.INIT_RAM_2A = 256'hB800280419AC180C018DD18CFF4C5C00018D040D218CFF4C018D040D658CFF4C;
defparam sp_inst_7.INIT_RAM_2B = 256'h018D240DA18CFF4C018D240DE58CFF4C29AC2C0C018D758CFF2C0180618CFF4C;
defparam sp_inst_7.INIT_RAM_2C = 256'hFF2CCC00018D340DC18CFF4C018D340D058CFF4C29AC300C018D958CFF2C0400;
defparam sp_inst_7.INIT_RAM_2D = 256'h018DD58CFF0C9400018D140DE18CFF4C018D140D258CFF4C29AC3C0C018DB58C;
defparam sp_inst_7.INIT_RAM_2E = 256'h19AC1C0C018DB18CFF4C5C00018D140D018CFF4C018D140D458CFF4C81AC400C;
defparam sp_inst_7.INIT_RAM_2F = 256'h818CFF4C018D280DC58CFF4C29AC2C0C018D558CFF0C0180418CFF4CB0002C04;
defparam sp_inst_7.INIT_RAM_30 = 256'h018D2C0DA18CFF4C018D2C0DE58CFF4C29AC300C018D758CFF0C0400018D280D;
defparam sp_inst_7.INIT_RAM_31 = 256'hFF0C9400018D140DC18CFF4C018D140D058CFF4C29AC3C0C018D958CFF0CCC00;
defparam sp_inst_7.INIT_RAM_32 = 256'h018D918CFF4C5C00018D140DE18CFF4C018D140D258CFF4C81AC400C018DB58C;
defparam sp_inst_7.INIT_RAM_33 = 256'h040D958CFF4C25AC400C018D258CFF0C10000180218CFF4CA8001C0419AC200C;
defparam sp_inst_7.INIT_RAM_34 = 256'h0180918CFF4C4400300419AC240C018D018CFF4C0000018D040D518CFF4C018D;
defparam sp_inst_7.INIT_RAM_35 = 256'hFF4CA400018D180DC18CFF4C018D180D058CFF4CC9AC400C018D958CFF0CE400;
defparam sp_inst_7.INIT_RAM_36 = 256'hFF4C6DAC400C018D058CFF0CE8000180018CFF4CE000340419AC280C018D718C;
defparam sp_inst_7.INIT_RAM_37 = 256'hFF4C7C00440419AC2C0C018DE18CFF4C4800018D1C0D318CFF4C018D1C0D758C;
defparam sp_inst_7.INIT_RAM_38 = 256'hF000018D300DB18CFF4C018D300DF58CFF4C29AC340C018D858CFF0C0180718C;
defparam sp_inst_7.INIT_RAM_39 = 256'hC58CFF0CB800018D1C0DD18CFF4C018D1C0D158CFF4C29AC380C018DA58CFF0C;
defparam sp_inst_7.INIT_RAM_3A = 256'h300C018DA18CFF4C8000018D1C0DF18CFF4C018D1C0D358CFF4CA5AC400C018D;
defparam sp_inst_7.INIT_RAM_3B = 256'h018D1C0DA58CFF4C49AC400C018D358CFF0C0180218CFF4C0400AC0038041DAC;
defparam sp_inst_7.INIT_RAM_3C = 256'hFF0C0180A18CFF4C4800400419AC340C018D118CFF4C2400018D1C0D618CFF4C;
defparam sp_inst_7.INIT_RAM_3D = 256'h018DD58CFF0CCC00018D380DE18CFF4C018D380D258CFF4C29AC340C018DB58C;
defparam sp_inst_7.INIT_RAM_3E = 256'h81AC400C018DF58CFF0C9400018D180D018CFF4C018D180D458CFF4C29AC380C;
defparam sp_inst_7.INIT_RAM_3F = 256'h780038041DAC380C018DD18CFF4C5C00018D180D218CFF4C018D180D658CFF4C;

SP sp_inst_8 (
    .DO({sp_inst_8_dout_w[15:0],sp_inst_8_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_8}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_8.READ_MODE = 1'b0;
defparam sp_inst_8.WRITE_MODE = 2'b01;
defparam sp_inst_8.BIT_WIDTH = 16;
defparam sp_inst_8.BLK_SEL = 3'b001;
defparam sp_inst_8.RESET_MODE = "SYNC";
defparam sp_inst_8.INIT_RAM_00 = 256'h180D918CFF4C018D180DD58CFF4C25AC400C018D658CFF0C0180518CFF4C4800;
defparam sp_inst_8.INIT_RAM_01 = 256'h040D918CFF4C018D040DD58CFF4C140048042DAC3C0C018D418CFF4C0000018D;
defparam sp_inst_8.INIT_RAM_02 = 256'h9000018D080DB18CFF4C018D080DF58CFF4CB5AC400C018D858CFF0CD3FF018D;
defparam sp_inst_8.INIT_RAM_03 = 256'hFF4C29AC2C0C018D058CFF0C0180F18CFF4C9C004C0419AC400C018D618CFF4C;
defparam sp_inst_8.INIT_RAM_04 = 256'h480D958CFF4C29AC300C018D258CFF0C3800018D440D318CFF4C018D440D758C;
defparam sp_inst_8.INIT_RAM_05 = 256'hFF4C018D140DB58CFF4C29AC3C0C018D458CFF0C0000018D480D518CFF4C018D;
defparam sp_inst_8.INIT_RAM_06 = 256'h140D918CFF4C018D140DD58CFF4CB5AC400C018D658CFF0CC800018D140D718C;
defparam sp_inst_8.INIT_RAM_07 = 256'h400D918CFF4C018D400DD58CFF4C940054042DAC440C018D418CFF4C9000018D;
defparam sp_inst_8.INIT_RAM_08 = 256'h2000018D400DB18CFF4C018D400DF58CFF4C45AC400C018D858CFF0CC7FF018D;
defparam sp_inst_8.INIT_RAM_09 = 256'hFF4C29AC340C018D058CFF0C0180F18CFF4C1C00500419AC480C018D618CFF4C;
defparam sp_inst_8.INIT_RAM_0A = 256'h400D958CFF2C29AC380C018D258CFF0CC800018D4C0D318CFF4C018D4C0D758C;
defparam sp_inst_8.INIT_RAM_0B = 256'hFF2C018D400DB58CFF2C7DAC400C018D458CFF0C9000018D400D518CFF2C018D;
defparam sp_inst_8.INIT_RAM_0C = 256'h018D400DA58CFF2C13FF4C00380431AC4C0C018D218CFF2C5800018D400D718C;
defparam sp_inst_8.INIT_RAM_0D = 256'h400D918CFF2C018D400DD58CFF2C0DAC400C018D658CFF0C018D400D618CFF2C;
defparam sp_inst_8.INIT_RAM_0E = 256'h018D040DA58CFF2C1FFF018D040D398CFF0C33FF1980018C898CFF0CE800018D;
defparam sp_inst_8.INIT_RAM_0F = 256'h0000D7FF0000DFFF0000E7FF0000EFFF0000F7FF0000FFFF018D040D618CFF2C;
defparam sp_inst_8.INIT_RAM_10 = 256'h000097FF00009FFF0000A7FF0000AFFF0000B7FF0000BFFF0000C7FF0000CFFF;
defparam sp_inst_8.INIT_RAM_11 = 256'h6076706180635FFF000067FF00006FFF000077FF00007FFF000087FF00008FFF;
defparam sp_inst_8.INIT_RAM_12 = 256'h1407210800681BFF0180018C31ACA18C006C898D7DAC540DBACCBACC008C8076;
defparam sp_inst_8.INIT_RAM_13 = 256'h2BFF7804180534063BFF4004180520064BFF000418051C06DBFF780400054006;
defparam sp_inst_8.INIT_RAM_14 = 256'h5804080500C600660807F3FF280400053C061C07B7FF00001BFFB80418053806;
defparam sp_inst_8.INIT_RAM_15 = 256'hA0041005240610078BFF5804100560C600660807C7FFA004080518060C07B7FF;
defparam sp_inst_8.INIT_RAM_16 = 256'h200418052C0608076FFFA0041805E00608075FFF58041805C0C6006608079BFF;
defparam sp_inst_8.INIT_RAM_17 = 256'hE0C6006608072BFF18040005340608073FFF580400058C060C0703FF4C005BFF;
defparam sp_inst_8.INIT_RAM_18 = 256'h100500C600660807EFFFE00408058C0608070FFFA00408051806EFFF58040805;
defparam sp_inst_8.INIT_RAM_19 = 256'h180510C600660807AFFF200410058C060807C3FFA004100524060807B3FF5804;
defparam sp_inst_8.INIT_RAM_1A = 256'h0005580617FF60006FFF200418058C06080783FFA0041805E006080773FF5804;
defparam sp_inst_8.INIT_RAM_1B = 256'h00041805B80608072FFFE804000518060C0743FF680400058406080763FF2804;
defparam sp_inst_8.INIT_RAM_1C = 256'h100793FFDC00EBFF00041805B8060807FFFF5004000558061407C3FF0C001BFF;
defparam sp_inst_8.INIT_RAM_1D = 256'h9FFF0004000558060C0763FFAC00BBFF3C04080574060807CFFF3C0408053806;
defparam sp_inst_8.INIT_RAM_1E = 256'h540063FF00041805B806080777FF80040005640608078BFFC00400058C060C07;
defparam sp_inst_8.INIT_RAM_1F = 256'hCFFF180033FF7C040805800643FF3C0408057C0647FF3C040805380610070BFF;
defparam sp_inst_8.INIT_RAM_20 = 256'hDFFFE00400058C060807FFFFA00400051806B3FFFC000BFF80040805A8061007;
defparam sp_inst_8.INIT_RAM_21 = 256'h0807AFFF200408051806B3FFA0040805C0060807A3FF58040805B0C600660807;
defparam sp_inst_8.INIT_RAM_22 = 256'h1005C80673FF20041005180677FFA0041005CC06080767FF58041005D0C60066;
defparam sp_inst_8.INIT_RAM_23 = 256'h0807D3FF1C002BFFA0041805980608071BFF58041805B0C60066080763FF6004;
defparam sp_inst_8.INIT_RAM_24 = 256'h0807BFFF5804080520C600660807FBFF200400058C0608070FFFA00400052406;
defparam sp_inst_8.INIT_RAM_25 = 256'h08077FFF5804100530C600660807BBFF2004080564060807CFFFA0040805C006;
defparam sp_inst_8.INIT_RAM_26 = 256'h00C60066080777FFA0041005C8067BFF20041005640608078FFFA0041005CC06;
defparam sp_inst_8.INIT_RAM_27 = 256'h180623FFA0040005C0060807E7FF30003FFFA0041805980608072FFF58041805;
defparam sp_inst_8.INIT_RAM_28 = 256'hD400E3FF1004000564060807F7FF90040005C0060807BBFF04001FFF20040005;
defparam sp_inst_8.INIT_RAM_29 = 256'h78040805C00608075FFFA800B7FFE0040805CC060807D7FFA0040805D4068BFF;
defparam sp_inst_8.INIT_RAM_2A = 256'h5FFF8C040005CC06080723FF6C0087FF38040805800697FFF80408057C069BFF;
defparam sp_inst_8.INIT_RAM_2B = 256'h2BFFB0041805DC063BFF00041805D8064BFF4C040005C8065BFF0C0400051806;
defparam sp_inst_8.INIT_RAM_2C = 256'hEBFF64040805C806EFFFE40408056406080703FF64040805CC060807C7FF1000;
defparam sp_inst_8.INIT_RAM_2D = 256'h0807A3FF64040805E006080767FFB000CBFFB0041805DC06DBFF00041805D806;
defparam sp_inst_8.INIT_RAM_2E = 256'h5FFF200400058C06080773FFA0040005E006080737FF80008FFFE40408056C06;
defparam sp_inst_8.INIT_RAM_2F = 256'h1FFF20040805E006080733FFA0040805C006080723FF58040805B0C600660807;
defparam sp_inst_8.INIT_RAM_30 = 256'hDFFF20041005E0060807F3FFA0041005CC060807E3FF58041005C0C600660807;
defparam sp_inst_8.INIT_RAM_31 = 256'h9400A3FFA00418059806080793FF5804180590C600660807DBFFA0041005C806;
defparam sp_inst_8.INIT_RAM_32 = 256'hD8066FFF64040805C80673FFE4040805E006080787FF64040805CC0608074BFF;
defparam sp_inst_8.INIT_RAM_33 = 256'hE006080727FFA0040005C0060807EBFF34004FFFB0041805DC065FFF00041805;
defparam sp_inst_8.INIT_RAM_34 = 256'h8ACC008CB3FF807660767061806300208063607670610000000013FF20040005;
defparam sp_inst_8.INIT_RAM_35 = 256'h898CB2CC51CEFF2E018D31AC898CA1ADFF2DFD8CB2CC4400B2CC100CF1808ACC;
defparam sp_inst_8.INIT_RAM_36 = 256'h0C050186140740088ACC018D918CFF2C8ACDBC0CB2CCB2CCFD8CB2CC018D31CC;
defparam sp_inst_8.INIT_RAM_37 = 256'h00000000000000000000000000000000000000008400A2CC918C1C6C9FFFB404;
defparam sp_inst_8.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_39 = 256'h92CCD58C182C8BFF0BFF3C04759FA2CDFD8DA2CC000000000000000000000000;
defparam sp_inst_8.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000008400;
defparam sp_inst_8.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_3C = 256'h607670610000018D180DD18CFF2C018D180D158CFF2C759F92CDFD8D92CC0000;
defparam sp_inst_8.INIT_RAM_3D = 256'h058CB2CC018031AC898CB2CC91ADFF2D2800B2C0807660767061806300208063;
defparam sp_inst_8.INIT_RAM_3E = 256'h00000000000000000000000000008400A2CCD58C182C6BFFD58D100CB2CDB2CC;
defparam sp_inst_8.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_9 (
    .DO({sp_inst_9_dout_w[15:0],sp_inst_9_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_9}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_9.READ_MODE = 1'b0;
defparam sp_inst_9.WRITE_MODE = 2'b01;
defparam sp_inst_9.BIT_WIDTH = 16;
defparam sp_inst_9.BLK_SEL = 3'b001;
defparam sp_inst_9.RESET_MODE = "SYNC";
defparam sp_inst_9.INIT_RAM_00 = 256'h180D958CFF2C759FA2CDFD8DA2CC000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_01 = 256'h008C6FFFC076A076B061406300208063607670610000018D180D518CFF2C018D;
defparam sp_inst_9.INIT_RAM_02 = 256'h200489AC018C31CC898C72CC91CEFF2E8ACD618D100C72CD72C071808ACC8ACC;
defparam sp_inst_9.INIT_RAM_03 = 256'h0000000000000000000000000000000000008400B2CCE58C472C67FFC3FFB7FF;
defparam sp_inst_9.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_05 = 256'h472CFFFF240443FFC3FF759FB2CDFD8DB2CC0000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_06 = 256'h00000000000000000000000000000000000000000000000000008400A2CCE58C;
defparam sp_inst_9.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_08 = 256'hBC00018D040DB58CFF2C018D040DF18CFF2C759FA2CDFD8DA2CC000000000000;
defparam sp_inst_9.INIT_RAM_09 = 256'h000000000000000000000000000000000000840092CC918C1C6CB3FF33FF1804;
defparam sp_inst_9.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0B = 256'hB0610000000087FF1004759F92CDFD8D92CC0000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0C = 256'h280C018DE58CFEECAD80018C258CFEECA2C0C076A076B06140630020C063A076;
defparam sp_inst_9.INIT_RAM_0D = 256'hC58CFEEC018DB18CFF0C31AD280C018D018CFF0C818D0C0C018D118CFF0C218D;
defparam sp_inst_9.INIT_RAM_0E = 256'h418CFF0C018DB18CFF0C31AD018CF18CFF0C018D81CC00070980B1AE280C018D;
defparam sp_inst_9.INIT_RAM_0F = 256'h92CE6400B2CCFD8C018C918CFF0C92CC018C118CFF0C018D018CFF0C058D018C;
defparam sp_inst_9.INIT_RAM_10 = 256'h04074008B58C8D8CB2CC92CC000709A035CC280D92CE42CC000709A0B5CC280D;
defparam sp_inst_9.INIT_RAM_11 = 256'h000000000000840082CC298C02CC9D80B2CCB2CCFD8CB2CC17FF01840C0542C6;
defparam sp_inst_9.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_13 = 256'h82CDFD8D82CC0000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_14 = 256'hBBFF01840C0540C600460807958C8D8C31ACB2CC018DF18CFF0C4400B2C0759F;
defparam sp_inst_9.INIT_RAM_15 = 256'h018D31AC898CB2CC21ADFF0D4400B2C0B1AC018CE18CFF0CB2CDB2CC058CB2CC;
defparam sp_inst_9.INIT_RAM_16 = 256'h018DD58CFEECB98D100CB2CDB2CC058CB2CC1C00A2CC040C11AC018C618CFF0C;
defparam sp_inst_9.INIT_RAM_17 = 256'h0000000000000000840072CCE58C472C53FFAFFFA3FF2004A180A2CC79AC2C0C;
defparam sp_inst_9.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_19 = 256'h759F72CDFD8D72CC000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1A = 256'h00000000000000000000000000000000840062CCE58C472CEBFF24042FFFAFFF;
defparam sp_inst_9.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1C = 256'h018D040DA18CFF0C759F62CDFD8D62CC00000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1D = 256'h1C6C3BFF87FF07FF1804D4000180B18CFF0C0180218CFF0C018D040D658CFF0C;
defparam sp_inst_9.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000840052CC918C;
defparam sp_inst_9.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_20 = 256'hFEEC3FFF14040180818CFEEC0180F18CFEEC759F52CDFD8D52CC000000000000;
defparam sp_inst_9.INIT_RAM_21 = 256'h0807B58C8D8CB2CC3400B2C00180B18CFEEC0180218CFEEC61AC300C018DB58C;
defparam sp_inst_9.INIT_RAM_22 = 256'h1DAC400C018DF58CFEECC98D0C0CB2CDB2CC058CB2CC67FF01840C0500C60046;
defparam sp_inst_9.INIT_RAM_23 = 256'hFEECC076A076B06140630020C063A076B06100000180F18CFEEC0180618CFEEC;
defparam sp_inst_9.INIT_RAM_24 = 256'h018D918CFEEC818D0C0C018DA18CFEECCD8D280C018D758CFEEC7180018CB58C;
defparam sp_inst_9.INIT_RAM_25 = 256'h818CFEEC018D81CC00070980B1AE280C018D558CFEEC018D418CFEEC31AD280C;
defparam sp_inst_9.INIT_RAM_26 = 256'hA2CC018CA18CFEEC018D918CFEEC058D018CD18CFEEC018D418CFEEC31AD018C;
defparam sp_inst_9.INIT_RAM_27 = 256'h09A035CC280DA2CE6ECC000709A0B5CC280DA2CE6C00B2CCFD8C018C218CFEEC;
defparam sp_inst_9.INIT_RAM_28 = 256'hB2CCFD8CB2CC33FF01A40C050186040740086ECC018DB58C8D8CB2CCA2CC0007;
defparam sp_inst_9.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000840092CC518C05AC9580B2CC;
defparam sp_inst_9.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2B = 256'hFEECE5AC2C0C018D058CFEEC759F92CDFD8D92CC000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2C = 256'h918C1C6C018D140DC18CFF0C018D140D058CFF0C63FF2004E9AC5C0C018D718C;
defparam sp_inst_9.INIT_RAM_2D = 256'h00000000000000000000000000000000000000000000000000000000840082CC;
defparam sp_inst_9.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2F = 256'h7BFF1804D7FFEC000180918CFEEC0180018CFEEC759F82CDFD8D82CC00000000;
defparam sp_inst_9.INIT_RAM_30 = 256'h00000000000000000000000000000000000000000000840072CC918C1C6CFBFF;
defparam sp_inst_9.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_32 = 256'h200D918CFF0C018D200DD58CFF0C759F72CDFD8D72CC00000000000000000000;
defparam sp_inst_9.INIT_RAM_33 = 256'hFEEC0180A18CFEEC61AC300C018D358CFECC0180E18CFEEC0180518CFEEC018D;
defparam sp_inst_9.INIT_RAM_34 = 256'hB2CC058CB2CCC7FF01840C0580C600460807B58C8D8CB2CC3400B2C00180318C;
defparam sp_inst_9.INIT_RAM_35 = 256'hB06100000180718CFEEC0180E18CFEEC1DAC400C018D758CFECCC98D0C0CB2CD;
defparam sp_inst_9.INIT_RAM_36 = 256'h2D8D280C018DF58CFECC1580018C358CFECC80766076706180630020C063A076;
defparam sp_inst_9.INIT_RAM_37 = 256'h018DD58CFECC018DC18CFEEC31AD280C018D118CFEEC818D0C0C018D218CFEEC;
defparam sp_inst_9.INIT_RAM_38 = 256'h018C518CFEEC018DC18CFEEC31AD018C018CFEEC018D81CC00070980B1AE280C;
defparam sp_inst_9.INIT_RAM_39 = 256'h280DA2CE6C00B2CCFD8C018CA18CFEECA2CC018C218CFEEC018D118CFEEC058D;
defparam sp_inst_9.INIT_RAM_3A = 256'h40088ECC018DB58C8D8CB2CCA2CC000709A035CC280DA2CE8ECC000709A0B5CC;
defparam sp_inst_9.INIT_RAM_3B = 256'h100C55AC2C0C018D058CFECC9580B2CCB2CCFD8CB2CC93FF01A40C0501860407;
defparam sp_inst_9.INIT_RAM_3C = 256'hB2CC018D31CC898CB2CC31CEFF0E018D31AC898C81ADFF0DFD8CB2CC4400B2CC;
defparam sp_inst_9.INIT_RAM_3D = 256'h0180518CFEEC0180C18CFEEC018D518CFF0C018D218CFEECBC0CB2CCB2CCFD8C;
defparam sp_inst_9.INIT_RAM_3E = 256'h000000000000000000000000000000000000840092CC918C1C6CEFFF3C047BFF;
defparam sp_inst_9.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_10 (
    .DO({sp_inst_10_dout_w[15:0],sp_inst_10_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_10}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_10.READ_MODE = 1'b0;
defparam sp_inst_10.WRITE_MODE = 2'b01;
defparam sp_inst_10.BIT_WIDTH = 16;
defparam sp_inst_10.BLK_SEL = 3'b001;
defparam sp_inst_10.RESET_MODE = "SYNC";
defparam sp_inst_10.INIT_RAM_00 = 256'hFF0C018D1C0DB58CFF0C759F92CDFD8D92CC0000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_01 = 256'h3400B2C00180718CFEEC0180E18CFEEC61AC300C018D758CFECC018D1C0D718C;
defparam sp_inst_10.INIT_RAM_02 = 256'h0000C98D0C0CB2CDB2CC058CB2CC57FF01840C05C0C600460807B58C8D8CB2CC;
defparam sp_inst_10.INIT_RAM_03 = 256'hB2CC018031AC898CB2CC31ADFF0D2800B2C08076707680630020806360767061;
defparam sp_inst_10.INIT_RAM_04 = 256'h00000000000000000000000000008400A2CC918C1C6CD58D100CB2CDB2CC058C;
defparam sp_inst_10.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_06 = 256'h1C0D958CFF0C759FA2CDFD8DA2CC000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_07 = 256'h5005A0C60046407620763061C0630020806370760000018D1C0D518CFF0C018D;
defparam sp_inst_10.INIT_RAM_08 = 256'h407620763061C06300204063207630610000D7FF8184D60C04052FFF70840044;
defparam sp_inst_10.INIT_RAM_09 = 256'hC063002040632076306100008BFF8184D60C0805E3FF408400446405D0C60046;
defparam sp_inst_10.INIT_RAM_0A = 256'h2076306100003FFF8184D60C100597FF10840044780500C60046407620763061;
defparam sp_inst_10.INIT_RAM_0B = 256'hF3FF8184D60C20054BFFE08400448C0530C60046407620763061C06300204063;
defparam sp_inst_10.INIT_RAM_0C = 256'h4005FFFFB0840044A00560C60046407620763061C06300204063207630610000;
defparam sp_inst_10.INIT_RAM_0D = 256'h0044B40590C60046407620763061C06300204063207630610000A7FF8184D60C;
defparam sp_inst_10.INIT_RAM_0E = 256'h0046407620763061C063002040632076306100005BFF8184D60C8005B3FF8084;
defparam sp_inst_10.INIT_RAM_0F = 256'h3061C063002040632076306100000FFF8184D60C000567FF50840044C805C0C6;
defparam sp_inst_10.INIT_RAM_10 = 256'h4063207630610000C3FF8184D60C00051BFF20840044E005F0C6004640762076;
defparam sp_inst_10.INIT_RAM_11 = 256'h000077FF8184D60C0005CFFFF0840044F40520C60046407620763061C0630020;
defparam sp_inst_10.INIT_RAM_12 = 256'hD60C000583FFC08400240C0550C60046407620763061C0630020406320763061;
defparam sp_inst_10.INIT_RAM_13 = 256'h90840024240580C60046407620763061C063002040632076306100002BFF8184;
defparam sp_inst_10.INIT_RAM_14 = 256'hB0C60046407620763061C06300204063207630610000DFFF8184D60C000537FF;
defparam sp_inst_10.INIT_RAM_15 = 256'h20763061C0630020406320763061000093FF8184D60C0005EBFF608400243C05;
defparam sp_inst_10.INIT_RAM_16 = 256'h0020406320763061000047FF8184D60C00259FFF308400245005E0C600464076;
defparam sp_inst_10.INIT_RAM_17 = 256'h30610000FBFF8184D60C004553FF00840024640510C60046407620763061C063;
defparam sp_inst_10.INIT_RAM_18 = 256'h8184D60C008507FFD08400247C0540C60046407620763061C063002040632076;
defparam sp_inst_10.INIT_RAM_19 = 256'hBBFFA0840024940570C60046407620763061C06300204063207630610000AFFF;
defparam sp_inst_10.INIT_RAM_1A = 256'hB005A0C60046407620763061C0630020406320763061000063FF8184D60C0105;
defparam sp_inst_10.INIT_RAM_1B = 256'h407620763061C0630020406320763061000017FF8184D60C02056FFF70840024;
defparam sp_inst_10.INIT_RAM_1C = 256'hC06300204063207630610000CBFF8184D60C040523FF40840024C805D0C60046;
defparam sp_inst_10.INIT_RAM_1D = 256'h2076306100007FFF8184D60C0805D7FF10840024E00500C60046407620763061;
defparam sp_inst_10.INIT_RAM_1E = 256'h33FF8184D60C10058BFFE0840024F80530C60046407620763061C06300204063;
defparam sp_inst_10.INIT_RAM_1F = 256'h20053FFFB0840024100560C60046407620763061C06300204063207630610000;
defparam sp_inst_10.INIT_RAM_20 = 256'h0024240590C60046407620763061C06300204063207630610000E7FF8184D60C;
defparam sp_inst_10.INIT_RAM_21 = 256'h0026407620763061C063002040632076306100009BFF8184D60C4005F3FF8084;
defparam sp_inst_10.INIT_RAM_22 = 256'h3061C063002040632076306100004FFF8184D60C8005A7FF508400243805C0C6;
defparam sp_inst_10.INIT_RAM_23 = 256'h406320763061000003FF8184D60C00055BFF208400245005F0C6002640762076;
defparam sp_inst_10.INIT_RAM_24 = 256'h0000B7FF8184D60C00050FFFF0840024680520C60026407620763061C0630020;
defparam sp_inst_10.INIT_RAM_25 = 256'hD60C0005C3FFC0840024800550C60026407620763061C0630020406320763061;
defparam sp_inst_10.INIT_RAM_26 = 256'h90840024980580C60026407620763061C063002040632076306100006BFF8184;
defparam sp_inst_10.INIT_RAM_27 = 256'hB0C60026407620763061C063002040632076306100001FFF8184D60C000577FF;
defparam sp_inst_10.INIT_RAM_28 = 256'h20763061C06300204063207630610000D3FF8184D60C00052BFF60840024B005;
defparam sp_inst_10.INIT_RAM_29 = 256'h0020406320763061000087FF8184D60C0005DFFF30840024C805E0C600264076;
defparam sp_inst_10.INIT_RAM_2A = 256'h306100003BFF8184D60C000593FF00840024E40510C60026407620763061C063;
defparam sp_inst_10.INIT_RAM_2B = 256'h8184D60C000547FFD0840024FC0540C60026407620763061C063002040632076;
defparam sp_inst_10.INIT_RAM_2C = 256'hFBFFA0840024140570C60026407620763061C06300204063207630610000EFFF;
defparam sp_inst_10.INIT_RAM_2D = 256'h000DF18CD60C807660767061806300204063207630610000A3FF8184D60C0005;
defparam sp_inst_10.INIT_RAM_2E = 256'hA2CD92CC018C818CD60CA2CC318C818CD60C9FFF30840024C40560C60026018D;
defparam sp_inst_10.INIT_RAM_2F = 256'h31AC898CB2CCB1AD002D2180058CB1ACB2CCA2CD4000B2C00000A2CCB1AC92CC;
defparam sp_inst_10.INIT_RAM_30 = 256'h60767061806300208063607670610000BD8D7C0CB2CDB2CC058CB2CC0181018C;
defparam sp_inst_10.INIT_RAM_31 = 256'h80630020806360767061000037FFB2CC018C118CD60C018D020DF18CD60C8076;
defparam sp_inst_10.INIT_RAM_32 = 256'hB6CC3D8C818C018C118CD68CBACCFD8C818CC18C018C118CD68C807660767061;
defparam sp_inst_10.INIT_RAM_33 = 256'h60767061000047FFF08400240185BACC018D3C0D118CD68C018D040DF18CD60C;
defparam sp_inst_10.INIT_RAM_34 = 256'h806370760000BECC018C098CD18C018D080DF18CD60C80767076806300208063;
defparam sp_inst_10.INIT_RAM_35 = 256'hF18CD60C018E118CD60CB2CC7D8CCD8C018C118CD60C80766076706180630020;
defparam sp_inst_10.INIT_RAM_36 = 256'h7BFF408400240180018C31ACE18C002C898DB2CC718D400CB2CD018DB5CDF00D;
defparam sp_inst_10.INIT_RAM_37 = 256'h018DB5CDFDADFEED118CD60C018E118CD60C5FFF708400243C000180118CD60C;
defparam sp_inst_10.INIT_RAM_38 = 256'hBECCBECC018C158CD40C80766076706180630020806360767061000000000800;
defparam sp_inst_10.INIT_RAM_39 = 256'h018CD10C2D80118CBECCCFFFC084002473FF00041980008C37FF00042980058C;
defparam sp_inst_10.INIT_RAM_3A = 256'h0184B6CCB6CC018CD00C2D80218CBECC018D100D0D8CD40C13FF0184BACCBACC;
defparam sp_inst_10.INIT_RAM_3B = 256'h3061C06300208063607670610000018DFC0D0D8CD40C018D200D0D8CD40CDFFF;
defparam sp_inst_10.INIT_RAM_3C = 256'h1670167016701554002040632076306100000FFF23FFB08400243FFF40762076;
defparam sp_inst_10.INIT_RAM_3D = 256'h15F415F415F415F415F415F415F415F4156C1670167016701670167016701670;
defparam sp_inst_10.INIT_RAM_3E = 256'h16701670167016701670167016701670167016701670167016701670167015F4;
defparam sp_inst_10.INIT_RAM_3F = 256'h1670167016701670167016701670167016701670167016701670167016701670;

SP sp_inst_11 (
    .DO({sp_inst_11_dout_w[15:0],sp_inst_11_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_11}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_11.READ_MODE = 1'b0;
defparam sp_inst_11.WRITE_MODE = 2'b01;
defparam sp_inst_11.BIT_WIDTH = 16;
defparam sp_inst_11.BLK_SEL = 3'b001;
defparam sp_inst_11.RESET_MODE = "SYNC";
defparam sp_inst_11.INIT_RAM_00 = 256'h16701670167016701474140C14E4167016701670167016701670167016701670;
defparam sp_inst_11.INIT_RAM_01 = 256'h151C16701670143C167013E016701670151C14AC167016701670167016701670;
defparam sp_inst_11.INIT_RAM_02 = 256'h14002241004100000305502236000864122A2400147F000700002F0000000000;
defparam sp_inst_11.INIT_RAM_03 = 256'h107F18004541464942007F423E453E000810000000000808006000003E081408;
defparam sp_inst_11.INIT_RAM_04 = 256'h510108140000141400410800365600000000494936493600097130493C004545;
defparam sp_inst_11.INIT_RAM_05 = 256'h20007F417F087F00494101097F0049491C227F00414136497F0011123E513200;
defparam sp_inst_11.INIT_RAM_06 = 256'h01010100494946297F00514106097F0041417F107F000C0240407F001408013F;
defparam sp_inst_11.INIT_RAM_07 = 256'h4040040204004141552A5500417F4345610070086314630038401F201F004040;
defparam sp_inst_11.INIT_RAM_08 = 256'h40007D4478047F00A4A40201080054547F483800444438447F00545400040000;
defparam sp_inst_11.INIT_RAM_09 = 256'h20400400545408047C0024241824FC00444478047C001804004000002810007D;
defparam sp_inst_11.INIT_RAM_0A = 256'h0000000000000000000000001414444C4400A0A04428440030401C201C004040;
defparam sp_inst_11.INIT_RAM_0B = 256'h18E008F01E21180030087000043F3F0478C0C040000000000C10100000300000;
defparam sp_inst_11.INIT_RAM_0C = 256'h00E00200201800000418000000000000000016102719211E0070F000211E2100;
defparam sp_inst_11.INIT_RAM_0D = 256'h000000000000B080000000000101010100000000020102024080404000074000;
defparam sp_inst_11.INIT_RAM_0E = 256'h0000100010200F001008E0000001600060800000000030000000000001010100;
defparam sp_inst_11.INIT_RAM_0F = 256'h0888F8003F240700F81000001120180048883000212230008808700020202000;
defparam sp_inst_11.INIT_RAM_10 = 256'h1008E00022211C00880870000000000038C8380011200F001888E00011201900;
defparam sp_inst_11.INIT_RAM_11 = 256'h40404040100801001020000000000000000000000030000000C0000011220000;
defparam sp_inst_11.INIT_RAM_12 = 256'h00E000001423180710E830C00136000008087000020420008040080004040404;
defparam sp_inst_11.INIT_RAM_13 = 256'h08E8F80810203F201008F80810201807080830C011203F207088F80827023C20;
defparam sp_inst_11.INIT_RAM_14 = 256'h0808080021013F200800F8081E221807380830C000033F2008E8F80820233F20;
defparam sp_inst_11.INIT_RAM_15 = 256'hF8F8F80820203F200000F80838263F201828F808007F80C008F8000020202000;
defparam sp_inst_11.INIT_RAM_16 = 256'h100810E001013F200808F8081020100F100810E018073F200800F8083F003F20;
defparam sp_inst_11.INIT_RAM_17 = 256'h0800F808002000000808081822213800080870000C033F208888F8085038180F;
defparam sp_inst_11.INIT_RAM_18 = 256'h38C838082C033020688018083C073C03080008F8010E0000C800780820201F00;
defparam sp_inst_11.INIT_RAM_19 = 256'h00FE02003806000000000C0040400000020200002020382038C8081000200000;
defparam sp_inst_11.INIT_RAM_1A = 256'h80800000000000000000020080808080000000000000000002020000007F4000;
defparam sp_inst_11.INIT_RAM_1B = 256'h8080000010200E008880000020200E008080000011203F000080F80822221900;
defparam sp_inst_11.INIT_RAM_1C = 256'h0000800020003F208080F80893946B0080800000202020008888800022221F00;
defparam sp_inst_11.INIT_RAM_1D = 256'h808080802020200000000800302D3F208080F8087F80C0009898000020202000;
defparam sp_inst_11.INIT_RAM_1E = 256'h808000001120FF800080808020201F008080000020003F2080808080203F3F20;
defparam sp_inst_11.INIT_RAM_1F = 256'h80008080202000008080800024243300808000000020202080808080A0200E00;
defparam sp_inst_11.INIT_RAM_20 = 256'h80008080310E200080808000300C300F80008080060801008000808010201F00;
defparam sp_inst_11.INIT_RAM_21 = 256'h0080020000FF000000FF00003F0000007C800000212221008080800006188180;
defparam sp_inst_11.INIT_RAM_22 = 256'h0000CEEDCAD3B0DDCA2000002020204B20202020000000000202060000004000;
defparam sp_inst_11.INIT_RAM_23 = 256'hD6200000B5ABBBC9CCC6D6200000A7CABCCDB8D6BCC20000D6CABBC3F7C6ABB4;
defparam sp_inst_11.INIT_RAM_24 = 256'hC6CE20200000C9ABB5F7CCC6D6200000D2C2F1CFC6CE20200000BAABBBAACCC6;
defparam sp_inst_11.INIT_RAM_25 = 256'hACB3F2D0D8B50000B0A7B2CFD5D820200000CEB8B5F7CBD0C32000002020A5C6;
defparam sp_inst_11.INIT_RAM_26 = 256'hA7D0DECEF8C7BABB0000B0A7BFC6D6D5C7200000DCB0E5B0FDB320200000B6B7;
defparam sp_inst_11.INIT_RAM_27 = 256'h0000C5BAE6B4A7D02020000020F3B4E5B6B420200000EDB4485346B4B6200000;
defparam sp_inst_11.INIT_RAM_28 = 256'h202000002020E2BFB8D620200000CEEDC2B3B1C2BC200000CEEDC8DAC6E6BC20;
defparam sp_inst_11.INIT_RAM_29 = 256'h00005BCC5AF85A145960582044490000CED0C2CFC8D8B72000002020EDB4D8B5;
defparam sp_inst_11.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2B = 256'h0101FFFC0000000000000000000000000000000000000080C0C0808000000000;
defparam sp_inst_11.INIT_RAM_2C = 256'h0000FEFFFFFF0F0FFFFFFFFF00000000000000000000000000000000F0FE0301;
defparam sp_inst_11.INIT_RAM_2D = 256'h000000000000000000003F7FFFFFFFFF7F7F0700000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2F = 256'h7BAC7AA4799C793878D477CC773483D400000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_30 = 256'h002A2E332E322E318310824081C880C080487FE47F147EB07DE07D7C7D187CB4;
defparam sp_inst_11.INIT_RAM_31 = 256'h8A408A1089E488F8881887FC87C087688738870886B485C8851484B08D100020;
defparam sp_inst_11.INIT_RAM_32 = 256'h2E0A00003E2073256E756425656E20200A0D8CE08C808B948B648B048AA88A6C;
defparam sp_inst_11.INIT_RAM_33 = 256'h7830656E68434B3A49686F742D0A0D0A2E2E2E2E2E2E544E54462E2E2E2E2E2E;
defparam sp_inst_11.INIT_RAM_34 = 256'h2E432E2E2E2E2E2E2E0A0D0A2E2E2E2E2E2E4C495F542E2E2E2E2E2E2E0A000A;
defparam sp_inst_11.INIT_RAM_35 = 256'h54206F4300002E7472726E696165207269546C6168706550000D2E2E2E2E2E2E;
defparam sp_inst_11.INIT_RAM_36 = 256'hA490A444A3F8A3ACA360A314A2C8A27CA230A1E4000A747072656920656C7265;
defparam sp_inst_11.INIT_RAM_37 = 256'hA950A904A8B8A86CA820A7D4A788A73CA6F0A6A4A658A60CA5C0A574A528A4DC;
defparam sp_inst_11.INIT_RAM_38 = 256'hAE04AE04AE04AE04AE04AE04AE04AE04ADB4AE04AB18AACCAA80AA34A9E8A99C;
defparam sp_inst_11.INIT_RAM_39 = 256'h616F675F7865656C61687269616F675F7865ADD0AE04AE04AE04AE04AE04AE04;
defparam sp_inst_11.INIT_RAM_3A = 256'h7865656C61687269616F675F7865656C61687269616F675F7865656C61687269;
defparam sp_inst_11.INIT_RAM_3B = 256'h61687269616F675F7865656C61687269616F675F7865656C61687269616F675F;
defparam sp_inst_11.INIT_RAM_3C = 256'h626F675F7865656C61687269626F675F7865656C61687269616F675F7865656C;
defparam sp_inst_11.INIT_RAM_3D = 256'h7865656C61687269626F675F7865656C61687269626F675F7865656C61687269;
defparam sp_inst_11.INIT_RAM_3E = 256'h61687269626F675F7865656C61687269626F675F7865656C61687269626F675F;
defparam sp_inst_11.INIT_RAM_3F = 256'h636F675F7865656C61687269636F675F7865656C61687269626F675F7865656C;

SP sp_inst_12 (
    .DO({sp_inst_12_dout_w[15:0],sp_inst_12_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_12}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_12.READ_MODE = 1'b0;
defparam sp_inst_12.WRITE_MODE = 2'b01;
defparam sp_inst_12.BIT_WIDTH = 16;
defparam sp_inst_12.BLK_SEL = 3'b001;
defparam sp_inst_12.RESET_MODE = "SYNC";
defparam sp_inst_12.INIT_RAM_00 = 256'h7865656C61687269636F675F7865656C61687269636F675F7865656C61687269;
defparam sp_inst_12.INIT_RAM_01 = 256'h61687269636F675F7865656C61687269636F675F7865656C61687269636F675F;
defparam sp_inst_12.INIT_RAM_02 = 256'h646F675F7865656C61687269646F675F7865656C61687269636F675F7865656C;
defparam sp_inst_12.INIT_RAM_03 = 256'h7865656C61687269646F675F7865656C61687269646F675F7865656C61687269;
defparam sp_inst_12.INIT_RAM_04 = 256'h61687269646F675F7865656C61687269646F675F7865656C61687269646F675F;
defparam sp_inst_12.INIT_RAM_05 = 256'h03680344000C034C032C0000656C61687865656C61687269646F675F7865656C;
defparam sp_inst_12.INIT_RAM_06 = 256'h7E009252FF0082847F004A48CC0800004949494900007E427E00321E94100350;
defparam sp_inst_12.INIT_RAM_07 = 256'h09094909880844241424147F44407F8000000000FF00FE0202020000F8008284;
defparam sp_inst_12.INIT_RAM_08 = 256'h000F80126722C8A899A80030302046230202420B420000011121A62A00008849;
defparam sp_inst_12.INIT_RAM_09 = 256'h090A893F60801E2292222CF41020001002000000000040444444404040404040;
defparam sp_inst_12.INIT_RAM_0A = 256'h4242434102029444244404E48C104F20102011210101E628202C242410200909;
defparam sp_inst_12.INIT_RAM_0B = 256'h090A893F60801E2292222CF41020408808083F10010280FE82F2C444840400F8;
defparam sp_inst_12.INIT_RAM_0C = 256'h102C8890000020A08282400040404F20102011210101E628202C242410200909;
defparam sp_inst_12.INIT_RAM_0D = 256'h15150010000044547F5444004240404055555555404017155755575517008041;
defparam sp_inst_12.INIT_RAM_0E = 256'hFF12100082428086A252820010105C5040405020400040487F4850004040007F;
defparam sp_inst_12.INIT_RAM_0F = 256'h102011210101E628202C242410200909090A893F60801E2292222CF410201012;
defparam sp_inst_12.INIT_RAM_10 = 256'h0300103F20001611FF1090901010000080400718800008088888F80808084F20;
defparam sp_inst_12.INIT_RAM_11 = 256'hFF9200051909D008D15210086888007F15150010000044547F54440042404020;
defparam sp_inst_12.INIT_RAM_12 = 256'h4242434102029444244404E48C1080400300030C4080000000E0010000007F80;
defparam sp_inst_12.INIT_RAM_13 = 256'h090A893F60801E2292222CF41020408808083F10010280FE82F2C444840400F8;
defparam sp_inst_12.INIT_RAM_14 = 256'h0D030D11818100101010101040004F20102011210101E628202C242410200909;
defparam sp_inst_12.INIT_RAM_15 = 256'h214020106080C80AFF0888880000402116216710478010F017D8FE02FE008141;
defparam sp_inst_12.INIT_RAM_16 = 256'h2F1181800000E424FF24E40460803F40010E88083010F010FF10080808084126;
defparam sp_inst_12.INIT_RAM_17 = 256'h4A4A4A4A0000A22AA3A4AAA66488007F02020202608000FE2222222200008181;
defparam sp_inst_12.INIT_RAM_18 = 256'h10102040808000C05252525200004444444410106020FE929292848484040000;
defparam sp_inst_12.INIT_RAM_19 = 256'h404040407C0000FC4040404000005845404440204000807FC94900004040804F;
defparam sp_inst_12.INIT_RAM_1A = 256'h27242720000000FEF212F2020000504845485820400062A324A400004040FC40;
defparam sp_inst_12.INIT_RAM_1B = 256'h404240204000FC04000200004040402001064C8208101828C80F9C642404007F;
defparam sp_inst_12.INIT_RAM_1C = 256'h212100FF1F000808180F40FFF80040403F00071880804046C040C05840404344;
defparam sp_inst_12.INIT_RAM_1D = 256'h27242720000000FEF212F2020000504845485820400062A324A4000040407F21;
defparam sp_inst_12.INIT_RAM_1E = 256'h7F0080404080F808F8001010101009047F802100040412921E3210006010007F;
defparam sp_inst_12.INIT_RAM_1F = 256'h15150000040444547F5444006010101212FF12133040242424A6A42400007F20;
defparam sp_inst_12.INIT_RAM_20 = 256'h404040400000000082828282000031097F811127FF002010E3242086FE00007F;
defparam sp_inst_12.INIT_RAM_21 = 256'h4444444401018242220622420200818989894121418100004949494900007840;
defparam sp_inst_12.INIT_RAM_22 = 256'h08168092672208080E0908103020FF4949490001440442444848901010100000;
defparam sp_inst_12.INIT_RAM_23 = 256'h284B00004202A888E98820901010007F15150010000044547F54440042408040;
defparam sp_inst_12.INIT_RAM_24 = 256'h4949000144044244484890101010020202024202020200222222242400008047;
defparam sp_inst_12.INIT_RAM_25 = 256'h0300030C4080000000E00100000040220804481040408080929292928080FF49;
defparam sp_inst_12.INIT_RAM_26 = 256'h08168092672208080E0908103020FF4949490001440442444848901010108040;
defparam sp_inst_12.INIT_RAM_27 = 256'h010E88083010F010FF10080808084126214020106080C80AFF08888800008040;
defparam sp_inst_12.INIT_RAM_28 = 256'h16216710478010F017D8FE02FE0081410D030D11818100101010101040003F40;
defparam sp_inst_12.INIT_RAM_29 = 256'h0202020200002808A8A8A8AC182008080808081E8808E0809292929200004021;
defparam sp_inst_12.INIT_RAM_2A = 256'h090906010608E628202C22232424007F15150010000044547F5444004240001E;
defparam sp_inst_12.INIT_RAM_2B = 256'h04040404040402F292929292020200FE4242FE00204020222222242400007F89;
defparam sp_inst_12.INIT_RAM_2C = 256'h04040404000000F010101010000040301010281000001611909090004040047F;
defparam sp_inst_12.INIT_RAM_2D = 256'h000F800000016098808E800780000001460A222242408000545456540000000F;
defparam sp_inst_12.INIT_RAM_2E = 256'h4040481000000404040400004040475841583F44180820504C5080FEFA02007F;
defparam sp_inst_12.INIT_RAM_2F = 256'h0000000000000000000D04D204D204D204D204D248001B0000000001FFFF4141;
defparam sp_inst_12.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000101;
defparam sp_inst_12.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_13 (
    .DO({sp_inst_13_dout_w[15:0],sp_inst_13_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_13}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_13.READ_MODE = 1'b0;
defparam sp_inst_13.WRITE_MODE = 2'b01;
defparam sp_inst_13.BIT_WIDTH = 16;
defparam sp_inst_13.BLK_SEL = 3'b001;
defparam sp_inst_13.RESET_MODE = "SYNC";
defparam sp_inst_13.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_14 (
    .DO({sp_inst_14_dout_w[15:0],sp_inst_14_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_14}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_14.READ_MODE = 1'b0;
defparam sp_inst_14.WRITE_MODE = 2'b01;
defparam sp_inst_14.BIT_WIDTH = 16;
defparam sp_inst_14.BLK_SEL = 3'b001;
defparam sp_inst_14.RESET_MODE = "SYNC";
defparam sp_inst_14.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_15 (
    .DO({sp_inst_15_dout_w[15:0],sp_inst_15_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_15}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_15.READ_MODE = 1'b0;
defparam sp_inst_15.WRITE_MODE = 2'b01;
defparam sp_inst_15.BIT_WIDTH = 16;
defparam sp_inst_15.BLK_SEL = 3'b001;
defparam sp_inst_15.RESET_MODE = "SYNC";
defparam sp_inst_15.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_16 (
    .DO({sp_inst_16_dout_w[15:0],sp_inst_16_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_16}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_16.READ_MODE = 1'b0;
defparam sp_inst_16.WRITE_MODE = 2'b01;
defparam sp_inst_16.BIT_WIDTH = 16;
defparam sp_inst_16.BLK_SEL = 3'b001;
defparam sp_inst_16.RESET_MODE = "SYNC";
defparam sp_inst_16.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_17 (
    .DO({sp_inst_17_dout_w[15:0],sp_inst_17_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_17}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_17.READ_MODE = 1'b0;
defparam sp_inst_17.WRITE_MODE = 2'b01;
defparam sp_inst_17.BIT_WIDTH = 16;
defparam sp_inst_17.BLK_SEL = 3'b001;
defparam sp_inst_17.RESET_MODE = "SYNC";
defparam sp_inst_17.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_18 (
    .DO({sp_inst_18_dout_w[15:0],sp_inst_18_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_18}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_18.READ_MODE = 1'b0;
defparam sp_inst_18.WRITE_MODE = 2'b01;
defparam sp_inst_18.BIT_WIDTH = 16;
defparam sp_inst_18.BLK_SEL = 3'b001;
defparam sp_inst_18.RESET_MODE = "SYNC";
defparam sp_inst_18.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_19 (
    .DO({sp_inst_19_dout_w[15:0],sp_inst_19_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_19}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_19.READ_MODE = 1'b0;
defparam sp_inst_19.WRITE_MODE = 2'b01;
defparam sp_inst_19.BIT_WIDTH = 16;
defparam sp_inst_19.BLK_SEL = 3'b001;
defparam sp_inst_19.RESET_MODE = "SYNC";
defparam sp_inst_19.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_20 (
    .DO({sp_inst_20_dout_w[15:0],sp_inst_20_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_20}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_20.READ_MODE = 1'b0;
defparam sp_inst_20.WRITE_MODE = 2'b01;
defparam sp_inst_20.BIT_WIDTH = 16;
defparam sp_inst_20.BLK_SEL = 3'b001;
defparam sp_inst_20.RESET_MODE = "SYNC";
defparam sp_inst_20.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_21 (
    .DO({sp_inst_21_dout_w[15:0],sp_inst_21_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_21}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_21.READ_MODE = 1'b0;
defparam sp_inst_21.WRITE_MODE = 2'b01;
defparam sp_inst_21.BIT_WIDTH = 16;
defparam sp_inst_21.BLK_SEL = 3'b001;
defparam sp_inst_21.RESET_MODE = "SYNC";
defparam sp_inst_21.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_22 (
    .DO({sp_inst_22_dout_w[15:0],sp_inst_22_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_22}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_22.READ_MODE = 1'b0;
defparam sp_inst_22.WRITE_MODE = 2'b01;
defparam sp_inst_22.BIT_WIDTH = 16;
defparam sp_inst_22.BLK_SEL = 3'b001;
defparam sp_inst_22.RESET_MODE = "SYNC";
defparam sp_inst_22.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_23 (
    .DO({sp_inst_23_dout_w[15:0],sp_inst_23_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_23}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_23.READ_MODE = 1'b0;
defparam sp_inst_23.WRITE_MODE = 2'b01;
defparam sp_inst_23.BIT_WIDTH = 16;
defparam sp_inst_23.BLK_SEL = 3'b001;
defparam sp_inst_23.RESET_MODE = "SYNC";
defparam sp_inst_23.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_24 (
    .DO({sp_inst_24_dout_w[15:0],sp_inst_24_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_24}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_24.READ_MODE = 1'b0;
defparam sp_inst_24.WRITE_MODE = 2'b01;
defparam sp_inst_24.BIT_WIDTH = 16;
defparam sp_inst_24.BLK_SEL = 3'b001;
defparam sp_inst_24.RESET_MODE = "SYNC";
defparam sp_inst_24.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_25 (
    .DO({sp_inst_25_dout_w[15:0],sp_inst_25_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_25}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_25.READ_MODE = 1'b0;
defparam sp_inst_25.WRITE_MODE = 2'b01;
defparam sp_inst_25.BIT_WIDTH = 16;
defparam sp_inst_25.BLK_SEL = 3'b001;
defparam sp_inst_25.RESET_MODE = "SYNC";
defparam sp_inst_25.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_26 (
    .DO({sp_inst_26_dout_w[15:0],sp_inst_26_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_26}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_26.READ_MODE = 1'b0;
defparam sp_inst_26.WRITE_MODE = 2'b01;
defparam sp_inst_26.BIT_WIDTH = 16;
defparam sp_inst_26.BLK_SEL = 3'b001;
defparam sp_inst_26.RESET_MODE = "SYNC";
defparam sp_inst_26.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_27 (
    .DO({sp_inst_27_dout_w[15:0],sp_inst_27_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_27}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_27.READ_MODE = 1'b0;
defparam sp_inst_27.WRITE_MODE = 2'b01;
defparam sp_inst_27.BIT_WIDTH = 16;
defparam sp_inst_27.BLK_SEL = 3'b001;
defparam sp_inst_27.RESET_MODE = "SYNC";
defparam sp_inst_27.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_28 (
    .DO({sp_inst_28_dout_w[15:0],sp_inst_28_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_28}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_28.READ_MODE = 1'b0;
defparam sp_inst_28.WRITE_MODE = 2'b01;
defparam sp_inst_28.BIT_WIDTH = 16;
defparam sp_inst_28.BLK_SEL = 3'b001;
defparam sp_inst_28.RESET_MODE = "SYNC";
defparam sp_inst_28.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_29 (
    .DO({sp_inst_29_dout_w[15:0],sp_inst_29_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_29}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_29.READ_MODE = 1'b0;
defparam sp_inst_29.WRITE_MODE = 2'b01;
defparam sp_inst_29.BIT_WIDTH = 16;
defparam sp_inst_29.BLK_SEL = 3'b001;
defparam sp_inst_29.RESET_MODE = "SYNC";
defparam sp_inst_29.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_30 (
    .DO({sp_inst_30_dout_w[15:0],sp_inst_30_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_30}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_30.READ_MODE = 1'b0;
defparam sp_inst_30.WRITE_MODE = 2'b01;
defparam sp_inst_30.BIT_WIDTH = 16;
defparam sp_inst_30.BLK_SEL = 3'b001;
defparam sp_inst_30.RESET_MODE = "SYNC";
defparam sp_inst_30.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_31 (
    .DO({sp_inst_31_dout_w[15:0],sp_inst_31_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_31}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_31.READ_MODE = 1'b0;
defparam sp_inst_31.WRITE_MODE = 2'b01;
defparam sp_inst_31.BIT_WIDTH = 16;
defparam sp_inst_31.BLK_SEL = 3'b001;
defparam sp_inst_31.RESET_MODE = "SYNC";
defparam sp_inst_31.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_32 (
    .DO({sp_inst_32_dout_w[15:0],sp_inst_32_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_32.READ_MODE = 1'b0;
defparam sp_inst_32.WRITE_MODE = 2'b01;
defparam sp_inst_32.BIT_WIDTH = 16;
defparam sp_inst_32.BLK_SEL = 3'b001;
defparam sp_inst_32.RESET_MODE = "SYNC";
defparam sp_inst_32.INIT_RAM_00 = 256'h15005FFF001003AA150003801500028029800010288000100385143850000015;
defparam sp_inst_32.INIT_RAM_01 = 256'h03BF15FF040003BF140004000015040014385FFF028029805800038D15000380;
defparam sp_inst_32.INIT_RAM_02 = 256'h00000000000000004C0006484C00547403BD1500040003800406038814EC0406;
defparam sp_inst_32.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_33 (
    .DO({sp_inst_33_dout_w[15:0],sp_inst_33_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_1}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_33.READ_MODE = 1'b0;
defparam sp_inst_33.WRITE_MODE = 2'b01;
defparam sp_inst_33.BIT_WIDTH = 16;
defparam sp_inst_33.BLK_SEL = 3'b001;
defparam sp_inst_33.RESET_MODE = "SYNC";
defparam sp_inst_33.INIT_RAM_00 = 256'h29BE29BE29BE29BE29BE29BF29BF29BF29BF29BF29BF29BF29BF29BF15000400;
defparam sp_inst_33.INIT_RAM_01 = 256'h440003404400034044000340440003404000036E040029BE29BE29BE29BE29BE;
defparam sp_inst_33.INIT_RAM_02 = 256'h5000549E5000549A5000549C5000549C5000549B5000549B4400036044000342;
defparam sp_inst_33.INIT_RAM_03 = 256'h28BE28BE28BF28BF28BF28BF28BF28BF28BF28BF28BF15005000549D40000341;
defparam sp_inst_33.INIT_RAM_04 = 256'h293F001502802980298002BF0648040028BE28BE28BE28BE28BE28BE28BE28BE;
defparam sp_inst_33.INIT_RAM_05 = 256'h29BE29BE29BE02812981298102BE4C0002802880288003405405157F00152A3F;
defparam sp_inst_33.INIT_RAM_06 = 256'h28BE500029BF29BF28BE500057FF028029BF001128BE640028BE400028BE29BE;
defparam sp_inst_33.INIT_RAM_07 = 256'h28BF29BF002A5C00002128BF28BE293E001002BF28BF0000002A5C00002128BF;
defparam sp_inst_33.INIT_RAM_08 = 256'h600028BF28BF500029BF001500130013001228BF28BF28BE47FF28BF29BF0280;
defparam sp_inst_33.INIT_RAM_09 = 256'h500000670280006728BF6000028028BF29BF00155000283E001002BF02BF28BF;
defparam sp_inst_33.INIT_RAM_0A = 256'h0281288128810015001563FF28BF29BF02BF28BF57FE001500670281006728BF;
defparam sp_inst_33.INIT_RAM_0B = 256'h28BF57FE00152A3F57FE02805C000280283F500029BF02802980298002BF4C00;
defparam sp_inst_33.INIT_RAM_0C = 256'h2980298002BE4C000280288028800015001547FF283F293F2A0028BF29BF0280;
defparam sp_inst_33.INIT_RAM_0D = 256'h500329BF29BF28BF29BF02BF0280298029802980298029802980298029BF0281;
defparam sp_inst_33.INIT_RAM_0E = 256'h02BF2800001028BF028028BF29BF02805C020280283F293F2A00001028BF28BF;
defparam sp_inst_33.INIT_RAM_0F = 256'h28BF29BF028028BF57FE0015288028BF4C002880001002AD1C00004068020281;
defparam sp_inst_33.INIT_RAM_10 = 256'h28BF500229BF028028BF29BF028028BF57FD00150067288028BF500229BF0280;
defparam sp_inst_33.INIT_RAM_11 = 256'h0280288028BF500229BF028028BF29BF028028BF57FD001528BF028000152880;
defparam sp_inst_33.INIT_RAM_12 = 256'h28BF02800015288028BF500129BF028028BF29BF028028BF57FC001528BF0280;
defparam sp_inst_33.INIT_RAM_13 = 256'h57FC001528BF02800015288028BF500129BF028028BF29BF028028BF57FC0015;
defparam sp_inst_33.INIT_RAM_14 = 256'h028028BF57FC001528BF02800015288028BF500129BF028028BF29BF028028BF;
defparam sp_inst_33.INIT_RAM_15 = 256'h500029BF29BF028028BF500129BF028028BF57FB0280500129BF028028BF29BF;
defparam sp_inst_33.INIT_RAM_16 = 256'h028028BF29BF028028BF29BF001002BF2800001028BF028028BF001C028028BF;
defparam sp_inst_33.INIT_RAM_17 = 256'h28BF500029BF53FD67FF02802800001028BF028028BF67FD02802800001028BF;
defparam sp_inst_33.INIT_RAM_18 = 256'h28BF028028BF29BF028028BF29BF001002BF2800001028BF028028BF001C0280;
defparam sp_inst_33.INIT_RAM_19 = 256'h5000034057FA028053FD67FF02802800001028BF028028BF67FD028028000010;
defparam sp_inst_33.INIT_RAM_1A = 256'h47FC2800001028BF28BF29BF028028BF57FA00152A3F57FA02805C000280283F;
defparam sp_inst_33.INIT_RAM_1B = 256'h00672A0028BF0340293F001529BF0280298002BF4C0002812880288000150015;
defparam sp_inst_33.INIT_RAM_1C = 256'h02802880034004010280298002BF4C0002802880034029002A3F28BF43FF0340;
defparam sp_inst_33.INIT_RAM_1D = 256'h29800380157F0280298002BF4C00028028800340040103800280298002BF4C00;
defparam sp_inst_33.INIT_RAM_1E = 256'h28800340298002800380157F298003BA14000380157F2980039014000380157F;
defparam sp_inst_33.INIT_RAM_1F = 256'h001003BA1400002A5C0000200280001C03B228BF29BF0280298002BF4C000280;
defparam sp_inst_33.INIT_RAM_20 = 256'h006703402A3F157F293F00150280298002BF4C0002802880034029800380157F;
defparam sp_inst_33.INIT_RAM_21 = 256'h02802980298002BF4C00028028800340290000670340157F006700442A3F2900;
defparam sp_inst_33.INIT_RAM_22 = 256'h00672A00157F0340290000670381157F00672A00157F57FF00152A3F293F0015;
defparam sp_inst_33.INIT_RAM_23 = 256'h0280298002BF4C00028028802880034043FF034000672A00157F034043FF0340;
defparam sp_inst_33.INIT_RAM_24 = 256'h034029000067001402BF157F00672A00157F290000670380157F00672A00157F;
defparam sp_inst_33.INIT_RAM_25 = 256'h00672A00157F290000670380157F00672A00157F0280298002BF4C0002802880;
defparam sp_inst_33.INIT_RAM_26 = 256'h29BF28BF29BF29BF29BF0280298002BF4C00028028800340290000670380157F;
defparam sp_inst_33.INIT_RAM_27 = 256'h4C0002802880001528BF47FF29BF02BF28BF2900006728BF29BF028028BF5000;
defparam sp_inst_33.INIT_RAM_28 = 256'h28BF02802881157F440028BF29BF28BF6000028028BF29BF29BF0280298002BF;
defparam sp_inst_33.INIT_RAM_29 = 256'h29810015157F0015001728BF02802881157F500029810014157F001500140017;
defparam sp_inst_33.INIT_RAM_2A = 256'h29810014157F00150014001728BF02802881157F440028BF29BF02BF28BF5000;
defparam sp_inst_33.INIT_RAM_2B = 256'h298002BF4C0002802880034029810015157F0015001728BF02802881157F5000;
defparam sp_inst_33.INIT_RAM_2C = 256'h0014001728BF02802881157F440028BF29BF28BF6000028028BF29BF29BF0280;
defparam sp_inst_33.INIT_RAM_2D = 256'h28BF500029810015157F0015001728BF02802881157F500029810014157F0015;
defparam sp_inst_33.INIT_RAM_2E = 256'h157F500029810014157F00150014001728BF02802881157F440028BF29BF02BF;
defparam sp_inst_33.INIT_RAM_2F = 256'h29BF0280298002BF4C0002802880034029810015157F0015001728BF02802881;
defparam sp_inst_33.INIT_RAM_30 = 256'h02805C00001728BF02800014001728BF02802881157F29BF28BF6000028028BF;
defparam sp_inst_33.INIT_RAM_31 = 256'h5C00001728BF02800014001728BF02802881157F29BF02BF28BF500000155000;
defparam sp_inst_33.INIT_RAM_32 = 256'h0280288D1CC7293F001502802980298002BF4C00028028800015001550000280;
defparam sp_inst_33.INIT_RAM_33 = 256'h29BF29BF0280298002BF4C0002802880288003405457029A1CC700152A3F2900;
defparam sp_inst_33.INIT_RAM_34 = 256'h28BF034029BF0280298002BF4C00028028800340298028BF001528BF288028BF;
defparam sp_inst_33.INIT_RAM_35 = 256'h28BF2980039A140028BF29BF0280298002BF4C0002802880034047FF29BF02BF;
defparam sp_inst_33.INIT_RAM_36 = 256'h03A0140329BF29BF0280298002BF4C000280288003402900028028BF29000280;
defparam sp_inst_33.INIT_RAM_37 = 256'h004428BF2900006728BF157F29BF02BF004428BF29BF028029000280157F29BF;
defparam sp_inst_33.INIT_RAM_38 = 256'h4C0002802880034029000280157F40002A0028BF290002BE157F29000067157F;
defparam sp_inst_33.INIT_RAM_39 = 256'h02802880034029000281157F5000290002BE157F400028BF29BF0280298002BF;
defparam sp_inst_33.INIT_RAM_3A = 256'h28800340290002BE157F500029000281157F400028BF29BF0280298002BF4C00;
defparam sp_inst_33.INIT_RAM_3B = 256'h034029000280157F29002A3F157F5400293F001502802980298002BF4C000280;
defparam sp_inst_33.INIT_RAM_3C = 256'h2A3F293F2A00157F500029BF293F2A00157F0280298002BF4C00028028802880;
defparam sp_inst_33.INIT_RAM_3D = 256'h157F400003402A3F293F2A00157F0280298002BF4C0002802880034047FF0340;
defparam sp_inst_33.INIT_RAM_3E = 256'h02802880034029800396154A157F0280298002BF4C0002802880034029000280;
defparam sp_inst_33.INIT_RAM_3F = 256'h0280028057FA0280028057FA0280028057FA0280028002802980298002BF4C00;

SP sp_inst_34 (
    .DO({sp_inst_34_dout_w[15:0],sp_inst_34_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_2}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_34.READ_MODE = 1'b0;
defparam sp_inst_34.WRITE_MODE = 2'b01;
defparam sp_inst_34.BIT_WIDTH = 16;
defparam sp_inst_34.BLK_SEL = 3'b001;
defparam sp_inst_34.RESET_MODE = "SYNC";
defparam sp_inst_34.INIT_RAM_00 = 256'h57F90280028057F90280028057F90280028057F90280028057F90280028057FA;
defparam sp_inst_34.INIT_RAM_01 = 256'h001557F90280001557F90280001557F90280001557F90280028057F902800015;
defparam sp_inst_34.INIT_RAM_02 = 256'h0340034003400340034003400340034003400340500029BF03BF140057F90280;
defparam sp_inst_34.INIT_RAM_03 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_04 = 256'h57F90280028057F90280028047FF29BF02BF28BF034003400340034003400340;
defparam sp_inst_34.INIT_RAM_05 = 256'h034057F90280001557F90280028057F90280028057F90280028057F902800280;
defparam sp_inst_34.INIT_RAM_06 = 256'h0399140057FB001502BF57FB001502BF02802980298002BF4C00028028802880;
defparam sp_inst_34.INIT_RAM_07 = 256'h03400340034003400340034003400340034003400340034003400340500029BF;
defparam sp_inst_34.INIT_RAM_08 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_09 = 256'h57F402802980298002BF4C00028028802880034047FF29BF02BF28BF03400340;
defparam sp_inst_34.INIT_RAM_0A = 256'h034003400340034003400340034003400340034003400340500029BF03991400;
defparam sp_inst_34.INIT_RAM_0B = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_0C = 256'h2980298002BF4C00028028802880034047FF29BF02BF28BF0340034003400340;
defparam sp_inst_34.INIT_RAM_0D = 256'h543F541F541C543E02802980298002BF4C00028028802880034057F502800280;
defparam sp_inst_34.INIT_RAM_0E = 256'h28802880034057F70280001502802980298002BF4C000280288028800340542B;
defparam sp_inst_34.INIT_RAM_0F = 256'h298002BF4C00028028802880034057F70280028002802980298002BF4C000280;
defparam sp_inst_34.INIT_RAM_10 = 256'h0340034003400340034003400340500029BF0399140057F60280028002802980;
defparam sp_inst_34.INIT_RAM_11 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_12 = 256'h57F60280001547FF29BF02BF28BF034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_13 = 256'h034003400340034003400340034003400340034003400340500029BF03991400;
defparam sp_inst_34.INIT_RAM_14 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_15 = 256'h0340500029BF0399140057F50280028047FF29BF02BF28BF0340034003400340;
defparam sp_inst_34.INIT_RAM_16 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_17 = 256'h28BF034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_18 = 256'h028002802980298002BF4C00028028802880034057F40280001547FF29BF02BF;
defparam sp_inst_34.INIT_RAM_19 = 256'h0340034003400340034003400340034003400340500029BF0399140057F40280;
defparam sp_inst_34.INIT_RAM_1A = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_1B = 256'h28802880034057F40280001547FF29BF02BF28BF034003400340034003400340;
defparam sp_inst_34.INIT_RAM_1C = 256'h028057F30280028057F30280028057F30280028002802980298002BF4C000280;
defparam sp_inst_34.INIT_RAM_1D = 256'h500029BF03A3140057FF02822982298202BD4C00028028802880034057F30280;
defparam sp_inst_34.INIT_RAM_1E = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_1F = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_20 = 256'h0340500029BF03A314004401001557F3028057F20280001547FF29BF02BF28BF;
defparam sp_inst_34.INIT_RAM_21 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_22 = 256'h28BF034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_23 = 256'h0340034003400340500029BF03A3140043FF001557F30280034047FF29BF02BF;
defparam sp_inst_34.INIT_RAM_24 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_25 = 256'h47FF29BF02BF28BF034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_26 = 256'h034003400340034003400340500029BF03A314004401001557F2028050150280;
defparam sp_inst_34.INIT_RAM_27 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_28 = 256'h0280034047FF29BF02BF28BF0340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_29 = 256'h034003400340034003400340034003400340500029BF03A3140043FF001557F1;
defparam sp_inst_34.INIT_RAM_2A = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_2B = 256'h001557F002805014028047FF29BF02BF28BF0340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_2C = 256'h03400340034003400340034003400340034003400340500029BF03A314004401;
defparam sp_inst_34.INIT_RAM_2D = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_2E = 256'h03A3140043FF001557F00280034047FF29BF02BF28BF03400340034003400340;
defparam sp_inst_34.INIT_RAM_2F = 256'h03400340034003400340034003400340034003400340034003400340500029BF;
defparam sp_inst_34.INIT_RAM_30 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_31 = 256'h500029BF03A314004401001557EF02805012028047FF29BF02BF28BF03400340;
defparam sp_inst_34.INIT_RAM_32 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_33 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_34 = 256'h034003400340500029BF03A3140043FF001557EE0280034047FF29BF02BF28BF;
defparam sp_inst_34.INIT_RAM_35 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_36 = 256'h29BF02BF28BF0340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_37 = 256'h0340500029BF03A314004401001557EE028057ED0280001557F95011028047FF;
defparam sp_inst_34.INIT_RAM_38 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_39 = 256'h28BF034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_3A = 256'h0340034003400340500029BF03A3140043FF001557ED0280034047FF29BF02BF;
defparam sp_inst_34.INIT_RAM_3B = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_3C = 256'h47FF29BF02BF28BF034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_3D = 256'h034003400340034003400340500029BF03A314004401001557EC0280500F0280;
defparam sp_inst_34.INIT_RAM_3E = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_34.INIT_RAM_3F = 256'h0280034047FF29BF02BF28BF0340034003400340034003400340034003400340;

SP sp_inst_35 (
    .DO({sp_inst_35_dout_w[15:0],sp_inst_35_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_3}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_35.READ_MODE = 1'b0;
defparam sp_inst_35.WRITE_MODE = 2'b01;
defparam sp_inst_35.BIT_WIDTH = 16;
defparam sp_inst_35.BLK_SEL = 3'b001;
defparam sp_inst_35.RESET_MODE = "SYNC";
defparam sp_inst_35.INIT_RAM_00 = 256'h034003400340034003400340034003400340500029BE03A3140043FF001557EB;
defparam sp_inst_35.INIT_RAM_01 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_02 = 256'h001557EB0280500E028047FF29BE02BF28BE0340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_03 = 256'h03400340034003400340034003400340034003400340500029BE03A314004401;
defparam sp_inst_35.INIT_RAM_04 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_05 = 256'h03A3140043FF001557EA0280034047FF29BE02BF28BE03400340034003400340;
defparam sp_inst_35.INIT_RAM_06 = 256'h03400340034003400340034003400340034003400340034003400340500029BE;
defparam sp_inst_35.INIT_RAM_07 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_08 = 256'h500029BE03A314004401001557E90280500C028047FF29BE02BF28BE03400340;
defparam sp_inst_35.INIT_RAM_09 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_0A = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_0B = 256'h034003400340500029BE03A3140043FF001557E90280034047FF29BE02BF28BE;
defparam sp_inst_35.INIT_RAM_0C = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_0D = 256'h29BE02BF28BE0340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_0E = 256'h0340500029BE03A314004401001557E8028057E70280001557F3500B028047FF;
defparam sp_inst_35.INIT_RAM_0F = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_10 = 256'h28BE034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_11 = 256'h0340034003400340500029BE03A3140043FF001557E70280034047FF29BE02BF;
defparam sp_inst_35.INIT_RAM_12 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_13 = 256'h47FF29BE02BF28BE034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_14 = 256'h034003400340034003400340500029BE03A314004401001557E60280500A0280;
defparam sp_inst_35.INIT_RAM_15 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_16 = 256'h0280034047FF29BE02BF28BE0340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_17 = 256'h034003400340034003400340034003400340500029BE03A3140043FF001557E6;
defparam sp_inst_35.INIT_RAM_18 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_19 = 256'h001557E502805008028047FF29BE02BF28BE0340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_1A = 256'h03400340034003400340034003400340034003400340500029BE03A314004401;
defparam sp_inst_35.INIT_RAM_1B = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_1C = 256'h03A3140043FF001557E40280034047FF29BE02BF28BE03400340034003400340;
defparam sp_inst_35.INIT_RAM_1D = 256'h03400340034003400340034003400340034003400340034003400340500029BE;
defparam sp_inst_35.INIT_RAM_1E = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_1F = 256'h500029BE03A314004401001557E402805007028047FF29BE02BF28BE03400340;
defparam sp_inst_35.INIT_RAM_20 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_21 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_22 = 256'h034003400340500029BE03A3140043FF001557E30280034047FF29BE02BF28BE;
defparam sp_inst_35.INIT_RAM_23 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_24 = 256'h29BE02BF28BE0340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_25 = 256'h0340500029BE03A314004401001557E2028057E10280001557ED5005028047FF;
defparam sp_inst_35.INIT_RAM_26 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_27 = 256'h28BE034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_28 = 256'h0340034003400340500029BE03A3140043FF001557E10280034047FF29BE02BF;
defparam sp_inst_35.INIT_RAM_29 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_2A = 256'h47FF29BE02BF28BE034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_2B = 256'h034003400340034003400340500029BE03A314004401001557E1028050040280;
defparam sp_inst_35.INIT_RAM_2C = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_2D = 256'h0280034047FF29BE02BF28BE0340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_2E = 256'h034003400340034003400340034003400340500029BD03A3140043FF001557E0;
defparam sp_inst_35.INIT_RAM_2F = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_30 = 256'h001557DF02805002028047FF29BD02BF28BD0340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_31 = 256'h03400340034003400340034003400340034003400340500029BD03A314004401;
defparam sp_inst_35.INIT_RAM_32 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_33 = 256'h03A3140043FF001557DF0280034047FF29BD02BF28BD03400340034003400340;
defparam sp_inst_35.INIT_RAM_34 = 256'h03400340034003400340034003400340034003400340034003400340500029BD;
defparam sp_inst_35.INIT_RAM_35 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_36 = 256'h500029BD03A314004401001557DE02805001028047FF29BD02BF28BD03400340;
defparam sp_inst_35.INIT_RAM_37 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_38 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_39 = 256'h034003400340500029BD03A3140043FF001557DD0280034047FF29BD02BF28BD;
defparam sp_inst_35.INIT_RAM_3A = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_3B = 256'h29BD02BF28BD0340034003400340034003400340034003400340034003400340;
defparam sp_inst_35.INIT_RAM_3C = 256'h0280293F001502802980298002BF4C00028228822882001500155000028047FF;
defparam sp_inst_35.INIT_RAM_3D = 256'h034057DD028057DF028057DF57DF00152A3F57DF57DF001557DF57DF028157DF;
defparam sp_inst_35.INIT_RAM_3E = 256'h028157DF57DF028157DE0280293F001502802980298002BF4C00028028802880;
defparam sp_inst_35.INIT_RAM_3F = 256'h02BF4C00028028802880034057DD028057DE028057DF57DE00152A3F57DF57DF;

SP sp_inst_36 (
    .DO({sp_inst_36_dout_w[15:0],sp_inst_36_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_4}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_36.READ_MODE = 1'b0;
defparam sp_inst_36.WRITE_MODE = 2'b01;
defparam sp_inst_36.BIT_WIDTH = 16;
defparam sp_inst_36.BLK_SEL = 3'b001;
defparam sp_inst_36.RESET_MODE = "SYNC";
defparam sp_inst_36.INIT_RAM_00 = 256'h034003400340034003400340034003400340500029BF03991400028029802980;
defparam sp_inst_36.INIT_RAM_01 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_36.INIT_RAM_02 = 256'h028057FE028057FE028247FF29BF02BF28BF0340034003400340034003400340;
defparam sp_inst_36.INIT_RAM_03 = 256'h028257FE028357FE028257FE028157FE028057FE001557FE028357FE028257FE;
defparam sp_inst_36.INIT_RAM_04 = 256'h028357FD028357FD001557FD028357FE028257FE028057FE028257FE028257FE;
defparam sp_inst_36.INIT_RAM_05 = 256'h028057FD028257FD028057FD028357FD028057FD028357FD028057FD028357FD;
defparam sp_inst_36.INIT_RAM_06 = 256'h006728BF29BF29BF02802980298002BF4C00028028802880034057FD028257FD;
defparam sp_inst_36.INIT_RAM_07 = 256'h0340006728BF57FD001500670380006703400067004428BF57FD0015006702BE;
defparam sp_inst_36.INIT_RAM_08 = 256'h293F001502802980298002BF4C00028028802880034057FD0015006703800067;
defparam sp_inst_36.INIT_RAM_09 = 256'h00152A3F500029BF57FC028057FC001557FC0015006702BE006728BF500029BF;
defparam sp_inst_36.INIT_RAM_0A = 256'h2880288003406FFF028028BF29BF028028BF6FFF028128BF29BF028028BF57FD;
defparam sp_inst_36.INIT_RAM_0B = 256'h2980298002BF4C00028028802880034057FF001502802980298002BF4C000280;
defparam sp_inst_36.INIT_RAM_0C = 256'h28BF500158010280580002802A3F29BF29BF29BF293F001529BF29BF29BF0280;
defparam sp_inst_36.INIT_RAM_0D = 256'h29BF57FE28BF28BF29BF028028BF29BF6C00028128BF29BF02BF2A00001028BF;
defparam sp_inst_36.INIT_RAM_0E = 256'h28BF29BF028028BF57FB00152A00001028BF0010001C028028BF02B31C005000;
defparam sp_inst_36.INIT_RAM_0F = 256'h28BF28BF500147FF2A00001028BF28BF29BF028028BF29BF028028BF6FFF0280;
defparam sp_inst_36.INIT_RAM_10 = 256'h500029BF57FD28BF28BF29BF028028BF29BF6C00028128BF29BF02BF2A000010;
defparam sp_inst_36.INIT_RAM_11 = 256'h6FFF028028BF29BF028028BF57FB00152A00001002B91C00001028BF004028BF;
defparam sp_inst_36.INIT_RAM_12 = 256'h2A00001002B71C000280001028BF004028BF500029BF57FD28BF0015028028BF;
defparam sp_inst_36.INIT_RAM_13 = 256'h28BF28BF29BF028028BF29BF028028BF6FFF028028BF29BF028028BF57FA0015;
defparam sp_inst_36.INIT_RAM_14 = 256'h001529BF29BF02802980298002BF4C000280288028800340034047FE2A000010;
defparam sp_inst_36.INIT_RAM_15 = 256'h00152A00001028BF02AA1CC75000293F57FC28BF28BF29BF00402A3F293F293F;
defparam sp_inst_36.INIT_RAM_16 = 256'h293F57FB28BF0015028028BF6FFF02802A3F293F02802A3F29BF028028BF57FA;
defparam sp_inst_36.INIT_RAM_17 = 256'h02802A3F293F02802A3F29BF028028BF57F900152A00001028BF02A91CC75000;
defparam sp_inst_36.INIT_RAM_18 = 256'h500029BF29BF29BF29BF29BF02802980298002BF4C0002802880288003406FFF;
defparam sp_inst_36.INIT_RAM_19 = 256'h028028BF57FE001528BF001500670010006728BF006728BF001028BF004028BF;
defparam sp_inst_36.INIT_RAM_1A = 256'h29BF29BF29BF02812980298002BF4C0002802880288003406BFF28BF28BF29BF;
defparam sp_inst_36.INIT_RAM_1B = 256'h29BF28BF29BF0280004428BF500029BF004428BF4400034028BF29BF29BF29BF;
defparam sp_inst_36.INIT_RAM_1C = 256'h28BF57F800152A00001028BF29BF028028BF500029BF28BF57FA28BF28BF5000;
defparam sp_inst_36.INIT_RAM_1D = 256'h4C0002812880288003406BFF28BF28BF29BF028028BF6BFF28BF28BF29BF0280;
defparam sp_inst_36.INIT_RAM_1E = 256'h29BF02BF2A3F29BF29BF293F0015293F0015001529BF29BF02802980298002BF;
defparam sp_inst_36.INIT_RAM_1F = 256'h28BF500029BF57F928BF28BF5C0002802A3F29BF028028BF29BF6C00028128BF;
defparam sp_inst_36.INIT_RAM_20 = 256'h28BF6FFF028028BF29BF028028BF57F700152A00001002AA1C00001028BF0040;
defparam sp_inst_36.INIT_RAM_21 = 256'h00152A00001002A81C000280001028BF004028BF500029BF57F928BF00150280;
defparam sp_inst_36.INIT_RAM_22 = 256'h28BF029F1C00500029BF57F828BF28BF50006FFF028028BF29BF028028BF57F7;
defparam sp_inst_36.INIT_RAM_23 = 256'h288003406FFF028028BF29BF028028BF57F600152A00001028BF0010001C0280;
defparam sp_inst_36.INIT_RAM_24 = 256'h28BF29BF001C28BF28BF500029BF028029BF29BF0280298002BF4C0002802880;
defparam sp_inst_36.INIT_RAM_25 = 256'h001529BF29BF29BF02802980298002BF4C0002802880001528BF47FF29BF02BF;
defparam sp_inst_36.INIT_RAM_26 = 256'h28BF001557FF0280001502BF001128BF2A3F500129BF29BF293F0015293F0015;
defparam sp_inst_36.INIT_RAM_27 = 256'h28BF6C0028BF001502BF2A3F440028BF29BF002A5C0000210280002A5C000021;
defparam sp_inst_36.INIT_RAM_28 = 256'h500057FD001528BF028000152A3F001028BF001C28BF0015006700442A3F4400;
defparam sp_inst_36.INIT_RAM_29 = 256'h00152A3F00670280006728BF001028BF001C28BF0015006700442A3F29BF0280;
defparam sp_inst_36.INIT_RAM_2A = 256'h02BF4C0002802880288003406BFE28BF2A3F29BF028028BF57FC001528BF0015;
defparam sp_inst_36.INIT_RAM_2B = 256'h500029BF28BF29BF28BF500028BF4400280028BF29BF28BF29BF29BF02802980;
defparam sp_inst_36.INIT_RAM_2C = 256'h280028BF280028BF4000280028BF4000280028BF29BF028028BF29BF028028BF;
defparam sp_inst_36.INIT_RAM_2D = 256'h028028800015001547FF280028BF29BF028028BF500028BF4400280028BF5BFF;
defparam sp_inst_36.INIT_RAM_2E = 256'h034029002A3F157F43FF034000672A00157F0340293F00150280298002BF4C00;
defparam sp_inst_36.INIT_RAM_2F = 256'h57FF028057FF028357CD28901CC70015028602802980298002BF4C0002802880;
defparam sp_inst_36.INIT_RAM_30 = 256'h57FF001500670044288002B81CC702802980298002BF4C000280288028800340;
defparam sp_inst_36.INIT_RAM_31 = 256'h02B71CC757FF001500670044288002B81CC757FF001500670044288002B81CC7;
defparam sp_inst_36.INIT_RAM_32 = 256'h2A3F293F001502802980298002BF4C00028028802880034057FE001500672880;
defparam sp_inst_36.INIT_RAM_33 = 256'h00150067004828BF29BF02802980298002BF4C00028028802880034057FE0015;
defparam sp_inst_36.INIT_RAM_34 = 256'h293F001502802980298002BF4C00028028802880034057FE0015006728BF57FE;
defparam sp_inst_36.INIT_RAM_35 = 256'h00442A7F297F001502802980298002BF4C00028028802880034057FE00152A3F;
defparam sp_inst_36.INIT_RAM_36 = 256'h2980298002BF4C00028028802880034057FD001500672A7F57FD00150067006F;
defparam sp_inst_36.INIT_RAM_37 = 256'h001028BF02B11CC7500029BF57FE57FD2900028028881CC729BF039C14000280;
defparam sp_inst_36.INIT_RAM_38 = 256'h29BF43FF034000672A00157F034067FF028028BF29BF028028BF57FD00152A00;
defparam sp_inst_36.INIT_RAM_39 = 256'h157F500029000067001502BE157F00672A00157F440028BF29BF02BF28BF5000;
defparam sp_inst_36.INIT_RAM_3A = 256'h1CC700672A00157F50002900001028BF28851CC7440028BF43FF034000672A00;
defparam sp_inst_36.INIT_RAM_3B = 256'h2A0028841CC76FFF028028BF29BF028028BF29BF039414002900001028BF2885;
defparam sp_inst_36.INIT_RAM_3C = 256'h57FE5424028002802980298002BF4C0002802880288000150280500000154400;
defparam sp_inst_36.INIT_RAM_3D = 256'h293F02BF29BF2A7F297F001502812980298002BF4C0002802880288000150015;
defparam sp_inst_36.INIT_RAM_3E = 256'h02AA1CC7293F00670044288002AA1CC7293F00670044288002AB1CC7293F0280;
defparam sp_inst_36.INIT_RAM_3F = 256'h00672A00157F0340293F293F0280293F0067288002AA1CC7293F006700442880;

SP sp_inst_37 (
    .DO({sp_inst_37_dout_w[15:0],sp_inst_37_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_5}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_37.READ_MODE = 1'b0;
defparam sp_inst_37.WRITE_MODE = 2'b01;
defparam sp_inst_37.BIT_WIDTH = 16;
defparam sp_inst_37.BLK_SEL = 3'b001;
defparam sp_inst_37.RESET_MODE = "SYNC";
defparam sp_inst_37.INIT_RAM_00 = 256'h0067001502BE157F00672A00157F440028BF29BF02BF28BF500029BF43FF0340;
defparam sp_inst_37.INIT_RAM_01 = 256'h157F50002900001028BF28BE1CC7440028BF43FF034000672A00157F50002900;
defparam sp_inst_37.INIT_RAM_02 = 256'h29BF2A7F542300152A00001028BF28BD1CC72900001028BF28BE1CC700672A00;
defparam sp_inst_37.INIT_RAM_03 = 256'h500028BF400028BF29BF57F928BC1CC7001502BF6FFF028028BF29BF028028BF;
defparam sp_inst_37.INIT_RAM_04 = 256'h57FB028057FB028057FA57FA02802980298002BF4C0002812880288000150015;
defparam sp_inst_37.INIT_RAM_05 = 256'h293F2A0028BF400028BF29BF57FD039C140057FC00152A7F297F028057FB0280;
defparam sp_inst_37.INIT_RAM_06 = 256'h57FA293F001502802980298002BF4C0002802880288000152A3F293F02BF5000;
defparam sp_inst_37.INIT_RAM_07 = 256'h00152A7F297F0280006F2A3F57F900152A3F57FB028057FB028057FA028057FA;
defparam sp_inst_37.INIT_RAM_08 = 256'h288000152A3F293F02BF5000293F2A0028BF400028BF29BF57FD039C140057FB;
defparam sp_inst_37.INIT_RAM_09 = 256'h028057FA028057FA028057FA028057F957F902802980298002BF4C0002802880;
defparam sp_inst_37.INIT_RAM_0A = 256'h293F02BF5000293F2A0028BF400028BF29BF57FC039C140057FA00152A7F297F;
defparam sp_inst_37.INIT_RAM_0B = 256'h57F9028057F9028057F957F802802980298002BF4C0002802880288000152A3F;
defparam sp_inst_37.INIT_RAM_0C = 256'h293F2A0028BF400028BF29BF57FC039C140057FA00152A7F297F028057FA0280;
defparam sp_inst_37.INIT_RAM_0D = 256'h293F0015001502802980298002BF4C0002802880288000152A3F293F02BF5000;
defparam sp_inst_37.INIT_RAM_0E = 256'h006F00442A7F57F700152A3F57F9028057F9028057F9028057F857F8297F0015;
defparam sp_inst_37.INIT_RAM_0F = 256'h006F0010006F0067006F00442A7F006F2A3F57F7001500672A7F57F700150067;
defparam sp_inst_37.INIT_RAM_10 = 256'h400028BF29BF57FB039C140057F900152A7F297F0280006F0010006F00672A7F;
defparam sp_inst_37.INIT_RAM_11 = 256'h02802980298002BF4C0002802880288000152A3F293F02BF5000293F2A0028BF;
defparam sp_inst_37.INIT_RAM_12 = 256'h57FA039C140057F800152A7F297F028057F8028057F8028057F8028057F757F7;
defparam sp_inst_37.INIT_RAM_13 = 256'h02BF4C0002802880288000152A3F293F02BF5000293F2A0028BF400028BF29BF;
defparam sp_inst_37.INIT_RAM_14 = 256'h57F7028057F657F6297F0015297F0015293F29BF001500150015028029802980;
defparam sp_inst_37.INIT_RAM_15 = 256'h001500672A7F57F600150067006F00442A7F57F600152A3F57F7028057F70280;
defparam sp_inst_37.INIT_RAM_16 = 256'h006F00442A7F006F2A3F57F5001500672A7F57F500150067006F00442A7F57F6;
defparam sp_inst_37.INIT_RAM_17 = 256'h0010006F00672A7F006F0010006F00442A7F006F0010006F00672A7F006F0010;
defparam sp_inst_37.INIT_RAM_18 = 256'h28BF293F2A0028BF400028BF29BF57F9039C140057F700152A7F297F0280006F;
defparam sp_inst_37.INIT_RAM_19 = 256'h2A00028028BF294028BF006F0010006F2A00028028BF006F0040006F2A000280;
defparam sp_inst_37.INIT_RAM_1A = 256'h00152A3F293F02BF5000294028BF006F0010006F2A00028028BF006F0040006F;
defparam sp_inst_37.INIT_RAM_1B = 256'h57EF028002800280028057EB293F001502802980298002BF4C00028028802880;
defparam sp_inst_37.INIT_RAM_1C = 256'h0340034003400340034003400340500029BF03BF140057EF0280028002810280;
defparam sp_inst_37.INIT_RAM_1D = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_37.INIT_RAM_1E = 256'h28802880034047FF29BF02BF28BF034003400340034003400340034003400340;
defparam sp_inst_37.INIT_RAM_1F = 256'h2A3F580602802A3F293F02802A3F293F293F293F02802980298002BF4C000280;
defparam sp_inst_37.INIT_RAM_20 = 256'h03BF140057ED028002800280028057EA4C002880001002891C00004068050280;
defparam sp_inst_37.INIT_RAM_21 = 256'h03400340034003400340034003400340034003400340034003400340500029BF;
defparam sp_inst_37.INIT_RAM_22 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_37.INIT_RAM_23 = 256'h2A3F293F001557F8028044002A3F293F001557F847FF29BF02BF28BF03400340;
defparam sp_inst_37.INIT_RAM_24 = 256'h5004293F0280293F57EC028102800281028057ED028002800280028057E94400;
defparam sp_inst_37.INIT_RAM_25 = 256'h0281028057EC028002800280028057E9500457FD00152A3F500457FD00152A3F;
defparam sp_inst_37.INIT_RAM_26 = 256'h028057E944002A3F293F001557F8028044002A3F293F001557F757EC02810280;
defparam sp_inst_37.INIT_RAM_27 = 256'h57FC00152A3F5003293F0280293F57EC028102800281028057EC028002800280;
defparam sp_inst_37.INIT_RAM_28 = 256'h57EB028102800281028057EB028002800280028057E8500357FC00152A3F5003;
defparam sp_inst_37.INIT_RAM_29 = 256'h57EB028102800281028057EB028002800280028057E844002A3F293F001557F8;
defparam sp_inst_37.INIT_RAM_2A = 256'h028057E85002293F028057EB028002800281028057EB028002800280028057E8;
defparam sp_inst_37.INIT_RAM_2B = 256'h03BF14005002293F57FB00152A3F57EB028002800281028057EB028002800280;
defparam sp_inst_37.INIT_RAM_2C = 256'h03400340034003400340034003400340034003400340034003400340500029BF;
defparam sp_inst_37.INIT_RAM_2D = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_37.INIT_RAM_2E = 256'h2A3F293F5001293F028044002A3F293F001557F747FF29BF02BF28BF03400340;
defparam sp_inst_37.INIT_RAM_2F = 256'h2A3F40002A3F293F5C0002802A3F293F001557CB5000293F0280500157FB0015;
defparam sp_inst_37.INIT_RAM_30 = 256'h028002B81C000280293F02802A3F680002832A3F293F5C0002802A3F293F02BF;
defparam sp_inst_37.INIT_RAM_31 = 256'h0015006F2A3F293F5FFF02802A3F57ED028002800015028002802A3F57E60280;
defparam sp_inst_37.INIT_RAM_32 = 256'h028002B61C00028057E9028002800280028057E644002A3F293F001557F60280;
defparam sp_inst_37.INIT_RAM_33 = 256'h034003400340500029BF03BF140057EC028002800015028002802A3F57E60280;
defparam sp_inst_37.INIT_RAM_34 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_37.INIT_RAM_35 = 256'h29BF02BF28BF0340034003400340034003400340034003400340034003400340;
defparam sp_inst_37.INIT_RAM_36 = 256'h03400340034003400340500029BF03BF1400034057F900152A3F293F500047FF;
defparam sp_inst_37.INIT_RAM_37 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_37.INIT_RAM_38 = 256'h53F947FF29BF02BF28BF03400340034003400340034003400340034003400340;
defparam sp_inst_37.INIT_RAM_39 = 256'h57E7028002800280028057E4293F02802980298002BF4C000280288028800340;
defparam sp_inst_37.INIT_RAM_3A = 256'h2A3F293F001557F2028047FF2A3F580202802A3F293F02802A3F293F001557F2;
defparam sp_inst_37.INIT_RAM_3B = 256'h57C754035425028057E344012A3F293F001557F6028000150281001502BF4402;
defparam sp_inst_37.INIT_RAM_3C = 256'h034003400340034003400340034003400340034003400340500029BF03BE1400;
defparam sp_inst_37.INIT_RAM_3D = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_37.INIT_RAM_3E = 256'h500029BF03BE140054240280540357C647FF29BF02BF28BF0340034003400340;
defparam sp_inst_37.INIT_RAM_3F = 256'h0340034003400340034003400340034003400340034003400340034003400340;

SP sp_inst_38 (
    .DO({sp_inst_38_dout_w[15:0],sp_inst_38_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_6}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_38.READ_MODE = 1'b0;
defparam sp_inst_38.WRITE_MODE = 2'b01;
defparam sp_inst_38.BIT_WIDTH = 16;
defparam sp_inst_38.BLK_SEL = 3'b001;
defparam sp_inst_38.RESET_MODE = "SYNC";
defparam sp_inst_38.INIT_RAM_00 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_01 = 256'h034003400340500029BF03BF140057C35424028057E2500047FF29BF02BF28BF;
defparam sp_inst_38.INIT_RAM_02 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_03 = 256'h29BF02BF28BF0340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_04 = 256'h02BF4C000280288028800340034053FD57E4028002800280028057E1500047FF;
defparam sp_inst_38.INIT_RAM_05 = 256'h29BF03BF140057F500152A3F500057C244002A3F293F001557F3028029802980;
defparam sp_inst_38.INIT_RAM_06 = 256'h0340034003400340034003400340034003400340034003400340034003405000;
defparam sp_inst_38.INIT_RAM_07 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_08 = 256'h28BF29BF02802980298002BF4C00028028802880034047FF29BF02BF28BF0340;
defparam sp_inst_38.INIT_RAM_09 = 256'h028028802880034057FF001502802980298002BF4C00028028802880034057B5;
defparam sp_inst_38.INIT_RAM_0A = 256'h02802980298002BF4C00028028802880034057FF028102802980298002BF4C00;
defparam sp_inst_38.INIT_RAM_0B = 256'h0340500029BF0399140002802980298002BF4C00028028802880034057FF0015;
defparam sp_inst_38.INIT_RAM_0C = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_0D = 256'h28BF034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_0E = 256'h03400340034003400340034003400340500029BF03911400540547FF29BF02BF;
defparam sp_inst_38.INIT_RAM_0F = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_10 = 256'h29BF03911400540547FF29BF02BF28BF03400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_11 = 256'h0340034003400340034003400340034003400340034003400340034003405000;
defparam sp_inst_38.INIT_RAM_12 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_13 = 256'h034003400340034003400340500029BF03911400540847FF29BF02BF28BF0340;
defparam sp_inst_38.INIT_RAM_14 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_15 = 256'h0340540647FF29BF02BF28BF0340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_16 = 256'h00000341000000402A3F293F293F001502802980298002BF4C00028028802880;
defparam sp_inst_38.INIT_RAM_17 = 256'h157F034043FF034000672A00157F034029002A3F157F57B3293F0000001502BE;
defparam sp_inst_38.INIT_RAM_18 = 256'h034043FF034000672A00157F03402900157F293F2A00157F47FF034000672A00;
defparam sp_inst_38.INIT_RAM_19 = 256'h0340034003400340500029BF028057B2293F2A00157F47FF034000672A00157F;
defparam sp_inst_38.INIT_RAM_1A = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_1B = 256'h47FF29BF02BF28BF034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_1C = 256'h2A3F293F0015293F0015001502802980298002BF4C0002802880288000152A3F;
defparam sp_inst_38.INIT_RAM_1D = 256'h157F034043FF034000672A00157F034029002A3F157F57B1293F034100670040;
defparam sp_inst_38.INIT_RAM_1E = 256'h43FF034000672A00157F034029002A3F157F293F2A00157F47FF034000672A00;
defparam sp_inst_38.INIT_RAM_1F = 256'h034003400340500029BF028057B1293F2A00157F47FF034000672A00157F0340;
defparam sp_inst_38.INIT_RAM_20 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_21 = 256'h29BF02BF28BF0340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_22 = 256'h293F293F0015293F0015001502802980298002BF4C00028028802880034047FF;
defparam sp_inst_38.INIT_RAM_23 = 256'h2880034057FE001500152A3F0067000000152A3F283F293F001557FC00152A3F;
defparam sp_inst_38.INIT_RAM_24 = 256'h57FC00152A3F293F293F0015293F0015001502802980298002BF4C0002802880;
defparam sp_inst_38.INIT_RAM_25 = 256'h28802880034057FD001500152A3F0067000000142A3F00000014283F293F0015;
defparam sp_inst_38.INIT_RAM_26 = 256'h0340034003400340500029BF028B57B10280028002802980298002BF4C000280;
defparam sp_inst_38.INIT_RAM_27 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_28 = 256'h47FF29BF02BF28BF034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_29 = 256'h0340034003400340034003400340034003400340500029BF028B57B002800015;
defparam sp_inst_38.INIT_RAM_2A = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_2B = 256'h57FC0280028057B00280028047FF29BF02BF28BF034003400340034003400340;
defparam sp_inst_38.INIT_RAM_2C = 256'h0340034003400340034003400340034003400340034003400340500029BF028B;
defparam sp_inst_38.INIT_RAM_2D = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_2E = 256'h57FB0280001557FB0280028057FB0280028047FF29BF02BF28BF034003400340;
defparam sp_inst_38.INIT_RAM_2F = 256'h02BF4C000280288028800015001557FB0280028157FB0280028057FB02800282;
defparam sp_inst_38.INIT_RAM_30 = 256'h0340034003400340034003400340500029BF028E57FB02800281028029802980;
defparam sp_inst_38.INIT_RAM_31 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_32 = 256'h001557F8028047FF29BF02BF28BF034003400340034003400340034003400340;
defparam sp_inst_38.INIT_RAM_33 = 256'h4C000280288028800340293F001557F8028057FB02800280440003402A3F293F;
defparam sp_inst_38.INIT_RAM_34 = 256'h29802980298002BF4C00028028802880034057FB0280028002802980298002BF;
defparam sp_inst_38.INIT_RAM_35 = 256'h580002802A3F293F293F293F02BF293F0015293F29BF29BF001529BF00150280;
defparam sp_inst_38.INIT_RAM_36 = 256'h001502BE2A3F03405000293F0280293F02815000293F0280293F02805C000280;
defparam sp_inst_38.INIT_RAM_37 = 256'h28BF500029BF57FA0280028257F90280001557FB0280028257F9028000150067;
defparam sp_inst_38.INIT_RAM_38 = 256'h57F8028000152A3F63FF28BF2A3F29BF028028BF57F9028000152A00001028BF;
defparam sp_inst_38.INIT_RAM_39 = 256'h29BF02BF28BF293F001557F7028029BF03A2140057FA028002825C0002802A3F;
defparam sp_inst_38.INIT_RAM_3A = 256'h0280400128BF57FA0280028243FF006700142A3F2A3F440003402A3F400028BF;
defparam sp_inst_38.INIT_RAM_3B = 256'h5C0002802A3F293F02BF40000340006700142A3F2A3F293F44000340001557F6;
defparam sp_inst_38.INIT_RAM_3C = 256'h00102A3F004002BF2A3F40002A3F293F0340001557F60280293F001557F60280;
defparam sp_inst_38.INIT_RAM_3D = 256'h293F02806C0002802A3F293F028044002A3F298028BF00402A3F5000298028BF;
defparam sp_inst_38.INIT_RAM_3E = 256'h500063FF28BF2A3F29BF028028BF2900001557F50280001028BF28BF500029BF;
defparam sp_inst_38.INIT_RAM_3F = 256'h02BF4C0002802880288028800015283F57F70280001557F802800282293F02BF;

SP sp_inst_39 (
    .DO({sp_inst_39_dout_w[15:0],sp_inst_39_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_7}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_39.READ_MODE = 1'b0;
defparam sp_inst_39.WRITE_MODE = 2'b01;
defparam sp_inst_39.BIT_WIDTH = 16;
defparam sp_inst_39.BLK_SEL = 3'b001;
defparam sp_inst_39.RESET_MODE = "SYNC";
defparam sp_inst_39.INIT_RAM_00 = 256'h2A3F57F80280028057F60280028057F802800280293F29BF0015028129802980;
defparam sp_inst_39.INIT_RAM_01 = 256'h028028BF4400283F293F001557FC0280001502800015001502BF02BF02BF293F;
defparam sp_inst_39.INIT_RAM_02 = 256'h0281288028800015283F293F02BF500029002A3F028028BF290028BF2A3F5C00;
defparam sp_inst_39.INIT_RAM_03 = 256'h57F80280028257F60280001557F802800280293F29BF02812980298002BF4C00;
defparam sp_inst_39.INIT_RAM_04 = 256'h283F293F001557FC0280001502800015001502BF02BF02BF293F0280293F02BE;
defparam sp_inst_39.INIT_RAM_05 = 256'h2A3F2A3F001002BF2A3F29002A3F001002BF001028BF2A3F2A3F5000293F4400;
defparam sp_inst_39.INIT_RAM_06 = 256'h293F02BF58002A3F2A3F001002BF2A3F6FFF02802A3F293F02802A3F293F0015;
defparam sp_inst_39.INIT_RAM_07 = 256'h28B81CC7297F02802980298002BF4C000281288028800015283F57F602800282;
defparam sp_inst_39.INIT_RAM_08 = 256'h0280006F006700442A0028B71CC74400001557FE28B81CC74400001557FD0281;
defparam sp_inst_39.INIT_RAM_09 = 256'h4C0002802880288000152A7F297F0010006F0340006F2A0028B71CC7006F001C;
defparam sp_inst_39.INIT_RAM_0A = 256'h001528BF29BF500029BF02804000001428BF2880157F29BF29BF0280298002BF;
defparam sp_inst_39.INIT_RAM_0B = 256'h2A000380157F2980001528BF157F2880157F29BF0280298002BF4C0002802880;
defparam sp_inst_39.INIT_RAM_0C = 256'h029C1CC729BF0280298002BF4C000280288003402900006703800380157F0067;
defparam sp_inst_39.INIT_RAM_0D = 256'h157F29000067157F004428BF290002BE157F29BF02BF002A5C00002128BF2880;
defparam sp_inst_39.INIT_RAM_0E = 256'h0280298002BF4C0002802880034029000280157F290002BF157F2900006728BF;
defparam sp_inst_39.INIT_RAM_0F = 256'h02BF4C0002802880034029002A3F157F43FF034000672A00157F0340293F0015;
defparam sp_inst_39.INIT_RAM_10 = 256'h290000670340157F00672A00157F293F02806C0002802A3F293F001502802980;
defparam sp_inst_39.INIT_RAM_11 = 256'h4C0002802880034029000067157F00000015000000402A3F000000672A00157F;
defparam sp_inst_39.INIT_RAM_12 = 256'h0280288028BF29002A3F0010288028BF288028BF293F001529BF0280298002BF;
defparam sp_inst_39.INIT_RAM_13 = 256'h288028BF298028BF0280288028BF298028BF6000288028BF288028BF298028BF;
defparam sp_inst_39.INIT_RAM_14 = 256'h288028BF288028BF298028BF0280288028BF298028BF288028BF6400288028BF;
defparam sp_inst_39.INIT_RAM_15 = 256'h140057AD57AC57AC57AA02802980298002BF4C00028028800340298028BF6000;
defparam sp_inst_39.INIT_RAM_16 = 256'h0340034003400340034003400340034003400340500029BF03BF140057FD0384;
defparam sp_inst_39.INIT_RAM_17 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_39.INIT_RAM_18 = 256'h0340500029BF03BF140057AD47FF29BF02BF28BF034003400340034003400340;
defparam sp_inst_39.INIT_RAM_19 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_39.INIT_RAM_1A = 256'h28BF034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_39.INIT_RAM_1B = 256'h1CC70015001557B057AC290002B21CC75C0C0280001557A5028047FF29BF02BF;
defparam sp_inst_39.INIT_RAM_1C = 256'h2A00028D1CC74C002880001002931C000040680C02802A00028E1CC7290002B1;
defparam sp_inst_39.INIT_RAM_1D = 256'h29000280028C1CC75C0002802A0002B01CC72900028D1CC7540D02805C000280;
defparam sp_inst_39.INIT_RAM_1E = 256'h028B1CC729000280028B1CC75C0C02802A0002AF1CC7500C29000280028C1CC7;
defparam sp_inst_39.INIT_RAM_1F = 256'h2A0002AD1CC72900028A1CC7540C02805C0002802A00028B1CC7500C29000280;
defparam sp_inst_39.INIT_RAM_20 = 256'h5C0002802A0002AC1CC7500B29000280028A1CC729000280028A1CC75C000280;
defparam sp_inst_39.INIT_RAM_21 = 256'h02881CC75C0002802A0002AC1CC7500B2900028002891CC72900028002891CC7;
defparam sp_inst_39.INIT_RAM_22 = 256'h2900028002871CC75C0B02802A0002AB1CC7500B2900028002881CC729000280;
defparam sp_inst_39.INIT_RAM_23 = 256'h5417290002861CC7540B02805C0002802A0002871CC7500B2900028002871CC7;
defparam sp_inst_39.INIT_RAM_24 = 256'h02851CC7500A2900028002851CC72900028002861CC75C0A02802A0002A91CC7;
defparam sp_inst_39.INIT_RAM_25 = 256'h02841CC75C0A02802A0002A81CC75419290002851CC7540B02805C0002802A00;
defparam sp_inst_39.INIT_RAM_26 = 256'h02831CC7540A02805C0002802A0002831CC7500A2900028002841CC729000280;
defparam sp_inst_39.INIT_RAM_27 = 256'h1CC7500A2900028002821CC72900028002831CC75C0002802A0002A61CC72900;
defparam sp_inst_39.INIT_RAM_28 = 256'h2A0002A41CC750092900028002811CC72900028002821CC75C0002802A0002A5;
defparam sp_inst_39.INIT_RAM_29 = 256'h5C0902802A0002A31CC750092900028002811CC72900028002811CC75C000280;
defparam sp_inst_39.INIT_RAM_2A = 256'h540902805C0002802A0002BF1CC750092900028002801CC72900028002801CC7;
defparam sp_inst_39.INIT_RAM_2B = 256'h2900028002BE1CC72900028002BE1CC75C0002802A0002A21CC7290002BF1CC7;
defparam sp_inst_39.INIT_RAM_2C = 256'h1CC750082900028002BD1CC72900028002BE1CC75C0002802A0002A11CC75009;
defparam sp_inst_39.INIT_RAM_2D = 256'h2A00029F1CC750082900028002BC1CC72900028002BD1CC75C0002802A0002A0;
defparam sp_inst_39.INIT_RAM_2E = 256'h5C0002802A0002BB1CC750082900028002BC1CC72900028002BC1CC75C080280;
defparam sp_inst_39.INIT_RAM_2F = 256'h02BA1CC72900028002BA1CC75C0002802A00029E1CC7290002BB1CC754080280;
defparam sp_inst_39.INIT_RAM_30 = 256'h2900028002B91CC72900028002B91CC75C0002802A00029D1CC7500829000280;
defparam sp_inst_39.INIT_RAM_31 = 256'h1CC750072900028002B81CC72900028002B91CC75C0002802A00029C1CC75007;
defparam sp_inst_39.INIT_RAM_32 = 256'h2A0002B71CC750072900028002B71CC72900028002B81CC75C0702802A00029B;
defparam sp_inst_39.INIT_RAM_33 = 256'h028002B61CC75C0702802A00029A1CC7541C290002B71CC7540702805C000280;
defparam sp_inst_39.INIT_RAM_34 = 256'h290002B51CC7540702805C0002802A0002B61CC750072900028002B61CC72900;
defparam sp_inst_39.INIT_RAM_35 = 256'h1CC750062900028002B41CC72900028002B51CC75C0602802A0002981CC7540F;
defparam sp_inst_39.INIT_RAM_36 = 256'h1CC75C0602802A0002971CC7541F290002B41CC7540602805C0002802A0002B4;
defparam sp_inst_39.INIT_RAM_37 = 256'h1CC7540602805C0002802A0002B21CC750062900028002B31CC72900028002B3;
defparam sp_inst_39.INIT_RAM_38 = 256'h50052900028002B11CC72900028002B11CC75C0002802A0002951CC7290002B2;
defparam sp_inst_39.INIT_RAM_39 = 256'h02931CC750052900028002B01CC72900028002B11CC75C0002802A0002941CC7;
defparam sp_inst_39.INIT_RAM_3A = 256'h02802A0002AF1CC750052900028002AF1CC72900028002B01CC75C0502802A00;
defparam sp_inst_39.INIT_RAM_3B = 256'h2900028002AE1CC75C0502802A0002921CC7290002AF1CC75422540502805C00;
defparam sp_inst_39.INIT_RAM_3C = 256'h1CC7290002AD1CC7540502805C0002802A0002AE1CC750052900028002AE1CC7;
defparam sp_inst_39.INIT_RAM_3D = 256'h2A00028F1CC750042900028002AC1CC72900028002AD1CC75C0002802A000290;
defparam sp_inst_39.INIT_RAM_3E = 256'h5C0402802A00028E1CC750042900028002AC1CC72900028002AC1CC75C000280;
defparam sp_inst_39.INIT_RAM_3F = 256'h540402805C0002802A0002AA1CC750042900028002AB1CC72900028002AB1CC7;

SP sp_inst_40 (
    .DO({sp_inst_40_dout_w[15:0],sp_inst_40_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_8}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_40.READ_MODE = 1'b0;
defparam sp_inst_40.WRITE_MODE = 2'b01;
defparam sp_inst_40.BIT_WIDTH = 16;
defparam sp_inst_40.BLK_SEL = 3'b001;
defparam sp_inst_40.RESET_MODE = "SYNC";
defparam sp_inst_40.INIT_RAM_00 = 256'h028002A91CC72900028002A91CC75C0402802A00028D1CC7290002AA1CC7540F;
defparam sp_inst_40.INIT_RAM_01 = 256'h028002A81CC72900028002A81CC7540402805C0002802A0002A91CC750042900;
defparam sp_inst_40.INIT_RAM_02 = 256'h50032900028002A71CC72900028002A71CC75C0302802A00028B1CC757DD2900;
defparam sp_inst_40.INIT_RAM_03 = 256'h1CC75C0002802A00028A1CC7290002A61CC7540302805C0002802A0002A71CC7;
defparam sp_inst_40.INIT_RAM_04 = 256'h028002A51CC75C0002802A0002891CC750032900028002A61CC72900028002A6;
defparam sp_inst_40.INIT_RAM_05 = 256'h1CC72900028002A41CC75C0002802A0002881CC750032900028002A51CC72900;
defparam sp_inst_40.INIT_RAM_06 = 256'h028002A31CC72900028002A31CC75C0202802A0002871CC750022900028002A4;
defparam sp_inst_40.INIT_RAM_07 = 256'h028002A21CC72900028002A21CC7540202805C0002802A0002A31CC750022900;
defparam sp_inst_40.INIT_RAM_08 = 256'h50022900028002A11CC72900028002A11CC75C0202802A0002851CC757D52900;
defparam sp_inst_40.INIT_RAM_09 = 256'h1CC75C0002802A0002841CC7290002A01CC7540202805C0002802A0002A11CC7;
defparam sp_inst_40.INIT_RAM_0A = 256'h0280029F1CC75C0002802A0002831CC750012900028002A01CC72900028002A0;
defparam sp_inst_40.INIT_RAM_0B = 256'h1CC729000280029E1CC75C0102802A0002821CC7500129000280029F1CC72900;
defparam sp_inst_40.INIT_RAM_0C = 256'h29000280029D1CC757DE540102805C0002802A00029E1CC7500129000280029E;
defparam sp_inst_40.INIT_RAM_0D = 256'h0280029C1CC729000280029C1CC75C0102802A0002801CC729000280029D1CC7;
defparam sp_inst_40.INIT_RAM_0E = 256'h29000280029B1CC757A02900028002BF1CC757BF44002A0002BF1CC750002900;
defparam sp_inst_40.INIT_RAM_0F = 256'h034053F2034053F2034053F2034053F2034053F2034053F229000280029B1CC7;
defparam sp_inst_40.INIT_RAM_10 = 256'h034053F2034053F2034053F2034053F2034053F2034053F2034053F2034053F2;
defparam sp_inst_40.INIT_RAM_11 = 256'h2980298002BF53F2034053F2034053F2034053F2034053F2034053F2034053F2;
defparam sp_inst_40.INIT_RAM_12 = 256'h028002971C0057BE4C0028800010029E1C000040680802802A7F297F00150280;
defparam sp_inst_40.INIT_RAM_13 = 256'h57C002810280028057C002800280028057C000150280028057C1028000150281;
defparam sp_inst_40.INIT_RAM_14 = 256'h02800280029C1C00028057C0028000150280028057BD500857C0028102800280;
defparam sp_inst_40.INIT_RAM_15 = 256'h028002800280028057BD02800280029B1C00028057C0028002800280028057BD;
defparam sp_inst_40.INIT_RAM_16 = 256'h028102800280028057C0028002800280028057BD02800280029A1C00028057C0;
defparam sp_inst_40.INIT_RAM_17 = 256'h02981C00028057C0028100150280028057C0028000150280028057BD500757C0;
defparam sp_inst_40.INIT_RAM_18 = 256'h028002981C00028057BF028002800280028057BF02800280028057BC02800280;
defparam sp_inst_40.INIT_RAM_19 = 256'h028002971C00028057BF028102800280028057BF028002800280028057BC0280;
defparam sp_inst_40.INIT_RAM_1A = 256'h0015028057BC500657BF028102800280028057BF028002800280028057BC0280;
defparam sp_inst_40.INIT_RAM_1B = 256'h001502800280028057BF028000150280028057BF028000150280028057BE0280;
defparam sp_inst_40.INIT_RAM_1C = 256'h028057BB500557BE001502800280028057BE028000150280028057BB500657BF;
defparam sp_inst_40.INIT_RAM_1D = 256'h57BE001500150280028057BB500557BE028102800280028057BE028002800281;
defparam sp_inst_40.INIT_RAM_1E = 256'h500557BE001502800280028057BE028100150280028057BE0280001502800280;
defparam sp_inst_40.INIT_RAM_1F = 256'h57BA500557BD02810280028057BD02810280028057BE028002800281028057BB;
defparam sp_inst_40.INIT_RAM_20 = 256'h57BD028000150280028057BC02800015028057BA500457BE0280028002800280;
defparam sp_inst_40.INIT_RAM_21 = 256'h028057BC02810280028057BD028002800280028057BA02800280028F1C000280;
defparam sp_inst_40.INIT_RAM_22 = 256'h0280028057BC02810280028057BD028002800280028057BA02800280028E1C00;
defparam sp_inst_40.INIT_RAM_23 = 256'h028057B9500457BD028002800280028057BA02800280028D1C00028057BC0281;
defparam sp_inst_40.INIT_RAM_24 = 256'h028057B902800280028C1C00028057BC028100150280028057BD028000150280;
defparam sp_inst_40.INIT_RAM_25 = 256'h028057B902800280028B1C00028057BC028102800280028057BC028002800280;
defparam sp_inst_40.INIT_RAM_26 = 256'h028A1C00028057BB02810280028057BC028102800280028057BC028002800280;
defparam sp_inst_40.INIT_RAM_27 = 256'h028057BC028000150280028057B8500357BC028002800280028057B902800280;
defparam sp_inst_40.INIT_RAM_28 = 256'h500257BB028100150280028057BB028000150280028057B8500357BB02810015;
defparam sp_inst_40.INIT_RAM_29 = 256'h028002800280028057B8500257BB028002800280028057BA02800280028057B8;
defparam sp_inst_40.INIT_RAM_2A = 256'h57BB028000150280028057B8500257BA02810280028057BA02800280028057BB;
defparam sp_inst_40.INIT_RAM_2B = 256'h57BA02810280028057BA00150280028057BA02810015028057BA028100150280;
defparam sp_inst_40.INIT_RAM_2C = 256'h57B902810280028057BA028002800280028057BB028002800280028057B75002;
defparam sp_inst_40.INIT_RAM_2D = 256'h028057BA028002800280028057B7500157B902810280028057B9001502800280;
defparam sp_inst_40.INIT_RAM_2E = 256'h57BA028100150280028057BA028000150280028057B7500157BA028002800280;
defparam sp_inst_40.INIT_RAM_2F = 256'h57BA028102800280028057BA028002800280028057B70280028002811C000280;
defparam sp_inst_40.INIT_RAM_30 = 256'h57B9028102800280028057B9028002800280028057B60280028002801C000280;
defparam sp_inst_40.INIT_RAM_31 = 256'h500057B9028002800280028057B60280028002BF1C00028057B8028102800280;
defparam sp_inst_40.INIT_RAM_32 = 256'h028057B802810280028057B9028002800280028057B9028002800280028057B6;
defparam sp_inst_40.INIT_RAM_33 = 256'h0280028057B9028000150280028057B5500057B802810280028057B800150280;
defparam sp_inst_40.INIT_RAM_34 = 256'h297F001557E402802980298002BF4C000280288028800340034057B902810015;
defparam sp_inst_40.INIT_RAM_35 = 256'h004028BF02B41CC728800010004002B41CC702BF28BF500029BF028040012A7F;
defparam sp_inst_40.INIT_RAM_36 = 256'h02800015028002802A7F298002B31CC72A7F63FF28BF29BF02BF28BF29800010;
defparam sp_inst_40.INIT_RAM_37 = 256'h0340034003400340034003400340034003400340500029BF03BF140057BB0280;
defparam sp_inst_40.INIT_RAM_38 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_40.INIT_RAM_39 = 256'h29BF03B21400579557F6028047FF29BF02BF28BF034003400340034003400340;
defparam sp_inst_40.INIT_RAM_3A = 256'h0340034003400340034003400340034003400340034003400340034003405000;
defparam sp_inst_40.INIT_RAM_3B = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_40.INIT_RAM_3C = 256'h2880288003402900028002AD1CC72900028002AE1CC747FF29BF02BF28BF0340;
defparam sp_inst_40.INIT_RAM_3D = 256'h028028BF29800010004028BF02AC1CC7500029BF02802980298002BF4C000280;
defparam sp_inst_40.INIT_RAM_3E = 256'h0340034003400340034003400340500029BF03B2140057946FFF028028BF29BF;
defparam sp_inst_40.INIT_RAM_3F = 256'h0340034003400340034003400340034003400340034003400340034003400340;

SP sp_inst_41 (
    .DO({sp_inst_41_dout_w[15:0],sp_inst_41_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_9}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_41.READ_MODE = 1'b0;
defparam sp_inst_41.WRITE_MODE = 2'b01;
defparam sp_inst_41.BIT_WIDTH = 16;
defparam sp_inst_41.BLK_SEL = 3'b001;
defparam sp_inst_41.RESET_MODE = "SYNC";
defparam sp_inst_41.INIT_RAM_00 = 256'h028002A91CC747FF29BF02BF28BF034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_01 = 256'h001557E102802980298002BF4C0002802880288003402900028002A91CC72900;
defparam sp_inst_41.INIT_RAM_02 = 256'h02805C0128800010004028BF02A71CC72A7F6802028028BF29BF40022A7F297F;
defparam sp_inst_41.INIT_RAM_03 = 256'h034003400340034003400340034003400340500029BF03BE1400579557D157F3;
defparam sp_inst_41.INIT_RAM_04 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_05 = 256'h140057F2028057D1579447FF29BF02BF28BF0340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_06 = 256'h0340034003400340034003400340034003400340034003400340500029BF03BE;
defparam sp_inst_41.INIT_RAM_07 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_08 = 256'h50002900028002A11CC72900028002A11CC747FF29BF02BF28BF034003400340;
defparam sp_inst_41.INIT_RAM_09 = 256'h034003400340034003400340034003400340500029BF03BF1400579157F20280;
defparam sp_inst_41.INIT_RAM_0A = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_0B = 256'h28800340034057F1028047FF29BF02BF28BF0340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_0C = 256'h02802A0002801CC740052A0002811CC729BF02802980298002BF4C0002802880;
defparam sp_inst_41.INIT_RAM_0D = 256'h02BF1CC7298028B21CC7001C0280288028B31CC768000280288028B31CC76802;
defparam sp_inst_41.INIT_RAM_0E = 256'h28B11CC7298028B11CC70010288028B11CC700150067002A5C00002102802A00;
defparam sp_inst_41.INIT_RAM_0F = 256'h28BF500029BF02BF288028B01CC729BF288028B11CC7298028B11CC702802880;
defparam sp_inst_41.INIT_RAM_10 = 256'h028002800280004028BF29BF002A5C000021028028BF29BF002A5C0000210280;
defparam sp_inst_41.INIT_RAM_11 = 256'h034003400340500029BF03B3140067FF28BF29BF02BF28BF57B50015028028BF;
defparam sp_inst_41.INIT_RAM_12 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_13 = 256'h29BF02BF28BF0340034003400340034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_14 = 256'h57AD00150280029C1C00028002800040001128BF288028AB1CC7500029BF47FF;
defparam sp_inst_41.INIT_RAM_15 = 256'h28800010004028BF02941CC7500029BF6BFF288028AA1CC728BF29BF028028BF;
defparam sp_inst_41.INIT_RAM_16 = 256'h2A0002B61CC76FFF028028BF29BF028028BF500029BF02805C00288028AA1CC7;
defparam sp_inst_41.INIT_RAM_17 = 256'h0340034003400340500029BF03BE1400579057CC57EE0280400128BF5C020280;
defparam sp_inst_41.INIT_RAM_18 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_19 = 256'h47FF29BF02BF28BF034003400340034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_1A = 256'h03400340034003400340034003400340500029BF03BE140057ED028057CC578F;
defparam sp_inst_41.INIT_RAM_1B = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_1C = 256'h29000280028D1CC747FF29BF02BF28BF03400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_1D = 256'h140057CB578C57ED02805000298028A21CC7298028A31CC729000280028D1CC7;
defparam sp_inst_41.INIT_RAM_1E = 256'h0340034003400340034003400340034003400340034003400340500029BF03BF;
defparam sp_inst_41.INIT_RAM_1F = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_20 = 256'h1CC757EC02802980289F1CC72980289F1CC747FF29BF02BF28BF034003400340;
defparam sp_inst_41.INIT_RAM_21 = 256'h02800280004028BF500029BF2980289E1CC72980289F1CC75C0002802A0002AC;
defparam sp_inst_41.INIT_RAM_22 = 256'h5C0002802A0002AA1CC767FF028028BF29BF028028BF57AA00150280028F1C00;
defparam sp_inst_41.INIT_RAM_23 = 256'h1CC702802980298002BF4C0002802880288003402980289C1CC72980289D1CC7;
defparam sp_inst_41.INIT_RAM_24 = 256'h2880289B1CC7680002802880289B1CC7680102802A0002A91CC740042A0002A9;
defparam sp_inst_41.INIT_RAM_25 = 256'h289A1CC700150067002A5C00002102802A0002A81CC72980289B1CC7001C0280;
defparam sp_inst_41.INIT_RAM_26 = 256'h29BF288028991CC7298028991CC70280288028991CC72980289A1CC700102880;
defparam sp_inst_41.INIT_RAM_27 = 256'h5C000020028028BF293F002A5C000020028028BF500029BF02BF288028991CC7;
defparam sp_inst_41.INIT_RAM_28 = 256'h29BF02BF28BF57AF00150280001502800280283F00150280004028BF29BF002A;
defparam sp_inst_41.INIT_RAM_29 = 256'h0340034003400340034003400340034003400340500029BF03A6140067FF28BF;
defparam sp_inst_41.INIT_RAM_2A = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_2B = 256'h1CC75C0102802A0002A21CC747FF29BF02BF28BF034003400340034003400340;
defparam sp_inst_41.INIT_RAM_2C = 256'h03BF14002900028002BD1CC72900028002BE1CC757E902805C00029128802894;
defparam sp_inst_41.INIT_RAM_2D = 256'h03400340034003400340034003400340034003400340034003400340500029BF;
defparam sp_inst_41.INIT_RAM_2E = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_2F = 256'h57E8028057A65000298028901CC7298028911CC747FF29BF02BF28BF03400340;
defparam sp_inst_41.INIT_RAM_30 = 256'h03400340034003400340034003400340034003400340500029BF03BF14005787;
defparam sp_inst_41.INIT_RAM_31 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_41.INIT_RAM_32 = 256'h028002B71CC72900028002B71CC747FF29BF02BF28BF03400340034003400340;
defparam sp_inst_41.INIT_RAM_33 = 256'h1CC72980288C1CC75C0002802A00029A1CC72980288C1CC72980288D1CC72900;
defparam sp_inst_41.INIT_RAM_34 = 256'h29BF028028BF57A50015028002BC1C0002800280004028BF500029BF2980288C;
defparam sp_inst_41.INIT_RAM_35 = 256'h288003402980288A1CC72980288A1CC75C0002802A0002981CC767FF028028BF;
defparam sp_inst_41.INIT_RAM_36 = 256'h680102802A0002961CC740032A0002971CC702802980298002BF4C0002802880;
defparam sp_inst_41.INIT_RAM_37 = 256'h2A0002951CC7298028881CC7001C0280288028891CC768000280288028891CC7;
defparam sp_inst_41.INIT_RAM_38 = 256'h288028871CC7298028871CC70010288028881CC700150067002A5C0000210280;
defparam sp_inst_41.INIT_RAM_39 = 256'h028028BF500029BF02BF288028861CC729BF288028871CC7298028871CC70280;
defparam sp_inst_41.INIT_RAM_3A = 256'h0280283F00150280004028BF29BF002A5C000020028028BF293F002A5C000020;
defparam sp_inst_41.INIT_RAM_3B = 256'h02805C0102802A0002921CC767FF28BF29BF02BF28BF57AA0015028000150280;
defparam sp_inst_41.INIT_RAM_3C = 256'h28BF29800010004028BF02AD1CC728800010004002AD1CC702BF28BF500029BF;
defparam sp_inst_41.INIT_RAM_3D = 256'h298028821CC7298028821CC7298002AC1CC7288028831CC763FF28BF29BF02BF;
defparam sp_inst_41.INIT_RAM_3E = 256'h034003400340034003400340034003400340500029BF03BF140057E402805784;
defparam sp_inst_41.INIT_RAM_3F = 256'h0340034003400340034003400340034003400340034003400340034003400340;

SP sp_inst_42 (
    .DO({sp_inst_42_dout_w[15:0],sp_inst_42_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_10}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_42.READ_MODE = 1'b0;
defparam sp_inst_42.WRITE_MODE = 2'b01;
defparam sp_inst_42.BIT_WIDTH = 16;
defparam sp_inst_42.BLK_SEL = 3'b001;
defparam sp_inst_42.RESET_MODE = "SYNC";
defparam sp_inst_42.INIT_RAM_00 = 256'h1CC72900028002A91CC747FF29BF02BF28BF0340034003400340034003400340;
defparam sp_inst_42.INIT_RAM_01 = 256'h500029BF298028BE1CC7298028BE1CC75C0002802A00028C1CC72900028002A9;
defparam sp_inst_42.INIT_RAM_02 = 256'h034067FF028028BF29BF028028BF57A20015028002AE1C0002800280004028BF;
defparam sp_inst_42.INIT_RAM_03 = 256'h28BF29800010004028BF02A61CC7500029BF0280298002BF4C00028028802880;
defparam sp_inst_42.INIT_RAM_04 = 256'h0340034003400340034003400340500029BF03BF14006FFF028028BF29BF0280;
defparam sp_inst_42.INIT_RAM_05 = 256'h0340034003400340034003400340034003400340034003400340034003400340;
defparam sp_inst_42.INIT_RAM_06 = 256'h028002A31CC747FF29BF02BF28BF034003400340034003400340034003400340;
defparam sp_inst_42.INIT_RAM_07 = 256'h028002B11C0002802980298002BF4C000280288003402900028002A31CC72900;
defparam sp_inst_42.INIT_RAM_08 = 256'h02802980298002BF4C000280288028800340577A0380157F0280577102AA1C00;
defparam sp_inst_42.INIT_RAM_09 = 256'h02BF4C000280288028800340577A0380157F0280577002A91C00028002B01C00;
defparam sp_inst_42.INIT_RAM_0A = 256'h288028800340577A0380157F0280577002A81C00028002B01C00028029802980;
defparam sp_inst_42.INIT_RAM_0B = 256'h57790380157F0280577002A61C00028002AF1C0002802980298002BF4C000280;
defparam sp_inst_42.INIT_RAM_0C = 256'h0280576F02A51C00028002AE1C0002802980298002BF4C000280288028800340;
defparam sp_inst_42.INIT_RAM_0D = 256'h1C00028002AD1C0002802980298002BF4C00028028802880034057790380157F;
defparam sp_inst_42.INIT_RAM_0E = 256'h1C0002802980298002BF4C00028028802880034057790380157F0280576F02A4;
defparam sp_inst_42.INIT_RAM_0F = 256'h298002BF4C00028028802880034057790380157F0281576F02A31C00028002AC;
defparam sp_inst_42.INIT_RAM_10 = 256'h028028802880034057780380157F0282576F02A21C00028002AB1C0002802980;
defparam sp_inst_42.INIT_RAM_11 = 256'h034057780380157F0284576E02A01C00028002AB1C0002802980298002BF4C00;
defparam sp_inst_42.INIT_RAM_12 = 256'h157F0288576E029F1C00028102AA1C0002802980298002BF4C00028028802880;
defparam sp_inst_42.INIT_RAM_13 = 256'h029E1C00028102A91C0002802980298002BF4C00028028802880034057780380;
defparam sp_inst_42.INIT_RAM_14 = 256'h02A81C0002802980298002BF4C00028028802880034057770380157F0290576E;
defparam sp_inst_42.INIT_RAM_15 = 256'h2980298002BF4C00028028802880034057770380157F03A0576D029D1C000281;
defparam sp_inst_42.INIT_RAM_16 = 256'h4C00028028802880034057770380157F1400576D029C1C00028102A71C000280;
defparam sp_inst_42.INIT_RAM_17 = 256'h2880034057760380157F1400576D029B1C00028102A71C0002802980298002BF;
defparam sp_inst_42.INIT_RAM_18 = 256'h0380157F1400576D02991C00028102A61C0002802980298002BF4C0002802880;
defparam sp_inst_42.INIT_RAM_19 = 256'h576C02981C00028102A51C0002802980298002BF4C0002802880288003405776;
defparam sp_inst_42.INIT_RAM_1A = 256'h028102A41C0002802980298002BF4C00028028802880034057760380157F1400;
defparam sp_inst_42.INIT_RAM_1B = 256'h02802980298002BF4C00028028802880034057760380157F1400576C02971C00;
defparam sp_inst_42.INIT_RAM_1C = 256'h02BF4C00028028802880034057750380157F1400576C02961C00028102A31C00;
defparam sp_inst_42.INIT_RAM_1D = 256'h28802880034057750380157F1400576B02951C00028102A31C00028029802980;
defparam sp_inst_42.INIT_RAM_1E = 256'h57750380157F1400576B02931C00028102A21C0002802980298002BF4C000280;
defparam sp_inst_42.INIT_RAM_1F = 256'h1400576B02921C00028202A11C0002802980298002BF4C000280288028800340;
defparam sp_inst_42.INIT_RAM_20 = 256'h1C00028202A01C0002802980298002BF4C00028028802880034057740380157F;
defparam sp_inst_42.INIT_RAM_21 = 256'h1C0002802980298002BF4C00028028802880034057740380157F1400576A0291;
defparam sp_inst_42.INIT_RAM_22 = 256'h298002BF4C00028028802880034057740380157F1400576A02901C000282029F;
defparam sp_inst_42.INIT_RAM_23 = 256'h028028802880034057740380157F1401576A028F1C000282029E1C0002802980;
defparam sp_inst_42.INIT_RAM_24 = 256'h034057730380157F1402576A028D1C000282029E1C0002802980298002BF4C00;
defparam sp_inst_42.INIT_RAM_25 = 256'h157F14045769028C1C000282029D1C0002802980298002BF4C00028028802880;
defparam sp_inst_42.INIT_RAM_26 = 256'h028B1C000282029C1C0002802980298002BF4C00028028802880034057730380;
defparam sp_inst_42.INIT_RAM_27 = 256'h029B1C0002802980298002BF4C00028028802880034057730380157F14085769;
defparam sp_inst_42.INIT_RAM_28 = 256'h2980298002BF4C00028028802880034057720380157F14105769028A1C000282;
defparam sp_inst_42.INIT_RAM_29 = 256'h4C00028028802880034057720380157F1420576802891C000282029A1C000280;
defparam sp_inst_42.INIT_RAM_2A = 256'h2880034057720380157F1440576802881C000282029A1C0002802980298002BF;
defparam sp_inst_42.INIT_RAM_2B = 256'h0380157F1480576802861C00028202991C0002802980298002BF4C0002802880;
defparam sp_inst_42.INIT_RAM_2C = 256'h576702851C00028302981C0002802980298002BF4C0002802880288003405771;
defparam sp_inst_42.INIT_RAM_2D = 256'h14020380157F02802980298002BF4C00028028802880034057710380157F1500;
defparam sp_inst_42.INIT_RAM_2E = 256'h28BF29BF28800380157F29BF28800380157F576702841C00028302971C002980;
defparam sp_inst_42.INIT_RAM_2F = 256'h0010004028BF02861C0040000340001728BF28BF500029BF034029BF001428BF;
defparam sp_inst_42.INIT_RAM_30 = 256'h2980298002BF4C0002802880288003406FFF028028BF29BF028028BF4C002880;
defparam sp_inst_42.INIT_RAM_31 = 256'h02BF4C000280288028800340577329BF28800380157F298014000380157F0280;
defparam sp_inst_42.INIT_RAM_32 = 256'h293F0340006728800380157F297F037F006F004428800380157F028029802980;
defparam sp_inst_42.INIT_RAM_33 = 256'h288028800340576602BF1C0000152A7F298002800380157F298014000380157F;
defparam sp_inst_42.INIT_RAM_34 = 256'h028028800340293F2A000380157F298014000380157F0280298002BF4C000280;
defparam sp_inst_42.INIT_RAM_35 = 256'h0380157F28800380157F29BF0340004428800380157F02802980298002BF4C00;
defparam sp_inst_42.INIT_RAM_36 = 256'h576502BD1C004C002880001002811C00004028BF6800028028BF298000141401;
defparam sp_inst_42.INIT_RAM_37 = 256'h2980001403BF15FF0380157F28800380157F576502BD1C00500029800380157F;
defparam sp_inst_42.INIT_RAM_38 = 256'h2A3F293F2A000380157F02802980298002BF4C00028028802880034003405000;
defparam sp_inst_42.INIT_RAM_39 = 256'h2880157F400003402A3F576402BB1C0057C402844000001557C4028440000340;
defparam sp_inst_42.INIT_RAM_3A = 256'h00152A3F293F2880157F400003402A3F290002800380157F576E00152A3F293F;
defparam sp_inst_42.INIT_RAM_3B = 256'h298002BF4C000280288028800340290002BF0380157F290002800380157F576D;
defparam sp_inst_42.INIT_RAM_3C = 256'h1C001C001C001C004C0002802880288003405768576402B91C00576802802980;
defparam sp_inst_42.INIT_RAM_3D = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_42.INIT_RAM_3E = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_42.INIT_RAM_3F = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;

SP sp_inst_43 (
    .DO({sp_inst_43_dout_w[15:0],sp_inst_43_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_11}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_43.READ_MODE = 1'b0;
defparam sp_inst_43.WRITE_MODE = 2'b01;
defparam sp_inst_43.BIT_WIDTH = 16;
defparam sp_inst_43.BLK_SEL = 3'b001;
defparam sp_inst_43.RESET_MODE = "SYNC";
defparam sp_inst_43.INIT_RAM_00 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_43.INIT_RAM_01 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_43.INIT_RAM_02 = 256'h3E08001C0000221C000000005549231362007F2A147F14000007000000000000;
defparam sp_inst_43.INIT_RAM_03 = 256'h27001214314B2100516100400000495102042000606008080800A00008080800;
defparam sp_inst_43.INIT_RAM_04 = 256'h0609020022411414140022140000000036361E290600494903050100494A3945;
defparam sp_inst_43.INIT_RAM_05 = 256'h41400041000008087A493E00090941497F00414122413E0049497C127C005949;
defparam sp_inst_43.INIT_RAM_06 = 256'h3F007F013149460019095E213E0009093E413E0008047F027F00404041227F00;
defparam sp_inst_43.INIT_RAM_07 = 256'h404040000102007F0000552A0041000049510708070008143F403F0040203F40;
defparam sp_inst_43.INIT_RAM_08 = 256'h84800040000004087CA41800097E185438004444204438004448785420000201;
defparam sp_inst_43.INIT_RAM_09 = 256'h3C00443F205448000408FC181800242438443800040878047C007F4100447F00;
defparam sp_inst_43.INIT_RAM_0A = 256'h0000F80000000000000000001414141454647CA01C0010283C403C0040207C20;
defparam sp_inst_43.INIT_RAM_0B = 256'h000000F00000FF200000FC880004040400404078000000000006060C00003300;
defparam sp_inst_43.INIT_RAM_0C = 256'h00001804004007000002E000000000000000000E1021242300008808001E031C;
defparam sp_inst_43.INIT_RAM_0D = 256'h00000000000000700000000000011F010000F00000020F010040F08000001820;
defparam sp_inst_43.INIT_RAM_0E = 256'h0000F810000F201000E008100000061804180000000000300000000001010101;
defparam sp_inst_43.INIT_RAM_0F = 256'h0008880800242404000020C0000E202000308808003024280070080800003F20;
defparam sp_inst_43.INIT_RAM_10 = 256'h00E00810001C21220070088800003F0000080808000E201100008810000E2021;
defparam sp_inst_43.INIT_RAM_11 = 256'h0040404000200402000840800000608000008000000030000000C000000F2231;
defparam sp_inst_43.INIT_RAM_12 = 256'h000038C0000B242700E028C80000300000F00848000108100000201000040404;
defparam sp_inst_43.INIT_RAM_13 = 256'h00108888000F202000E008080008202000380808000E20200000888820380223;
defparam sp_inst_43.INIT_RAM_14 = 256'h0000F808203F012108F800080002202000000808000000200010888800182020;
defparam sp_inst_43.INIT_RAM_15 = 256'h000800F80030202000000008002001200008C088000080800008080800003F20;
defparam sp_inst_43.INIT_RAM_16 = 256'h00E008080000012100F00808000F202000E00808003F002008F8C03000203F00;
defparam sp_inst_43.INIT_RAM_17 = 256'h08F8000800003F200018F808001C2120003808882030002000708888004F2424;
defparam sp_inst_43.INIT_RAM_18 = 256'h000800C82030032C081880680003000700F8F8000000380708380088001F2020;
defparam sp_inst_43.INIT_RAM_19 = 256'h0000020200C001000000C03000407F000002FE00001821260008080800003F20;
defparam sp_inst_43.INIT_RAM_1A = 256'h0000808000000000000004028080808000000000000000000004020400004040;
defparam sp_inst_43.INIT_RAM_1B = 256'h00008080203F201100F880000011201100008000000E201100008000203F2224;
defparam sp_inst_43.INIT_RAM_1C = 256'h00009898203F002100008000006094940080808000003F201888F08000132222;
defparam sp_inst_43.INIT_RAM_1D = 256'h0080808000003F200000F8080020022400800000000080800000800000003F20;
defparam sp_inst_43.INIT_RAM_1E = 256'h00808000000E20A100008000001F202000008080203F0021000080003F000020;
defparam sp_inst_43.INIT_RAM_1F = 256'h0080000000001F000000E08000192424008080800001213F0080008080FF2011;
defparam sp_inst_43.INIT_RAM_20 = 256'h8080008000202E3100800080000F030C808080000001300E80800080203F2020;
defparam sp_inst_43.INIT_RAM_21 = 256'h00007C020000000000000000404000000202000000302C30008080800001708E;
defparam sp_inst_43.INIT_RAM_22 = 256'h000020F3B4D5BDFCBEFD0000202020204F202020000000000404010100003F40;
defparam sp_inst_43.INIT_RAM_23 = 256'hCEB8000020ADCCF2B8ABCEB80000DCB0F1CFC6CEEBC80000B8D6D0D3CFC9D0B8;
defparam sp_inst_43.INIT_RAM_24 = 256'hBBB2B8D6000020D9CCE3D5D8CEB800002020ABCCBCCDB8D6000020FDCCF2CAAB;
defparam sp_inst_43.INIT_RAM_25 = 256'hF6B3C5BAB7D6000020DCCAA2BAF7CC20000020C6D6BDCBD1D3BB00002020E4C5;
defparam sp_inst_43.INIT_RAM_26 = 256'hBCCDD0D3DAC4E5B3000020DCCAE2CEB8BFE500002020A7CAA3C4BEC90000A7CE;
defparam sp_inst_43.INIT_RAM_27 = 256'h00002020F7C6C4BCDECE00002020CEEDD2A8CE2000002020F6B3414CD0C10000;
defparam sp_inst_43.INIT_RAM_28 = 256'h202000002020FAC2C6CE2020000020F3B4EBD2BECAC7000020F3B4DDC4F7B4C4;
defparam sp_inst_43.INIT_RAM_29 = 256'h00001C001C001C001C001C00003A000020F3D3EBC8B7BBB500002020F3CEB7D6;
defparam sp_inst_43.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_2B = 256'h01000307000000000000000000000000000000000000000080C0C0C000000000;
defparam sp_inst_43.INIT_RAM_2C = 256'h00000000FFFFFF9F0F9FFFFFFE0000000000000000000000000000000000FF07;
defparam sp_inst_43.INIT_RAM_2D = 256'h00000000000000000000071F7FFFF8F8FFFF3F1F000000000000000000000000;
defparam sp_inst_43.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_2F = 256'h1C001C001C001C001C001C001C001C0000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_30 = 256'h00000000000000001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_43.INIT_RAM_31 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C000000;
defparam sp_inst_43.INIT_RAM_32 = 256'h2E2E00000A0D20203A636620203A696C3C201C001C001C001C001C001C001C00;
defparam sp_inst_43.INIT_RAM_33 = 256'h78253A6C6E617965746E63752D2D00002E2E2E2E2E2E2E2E495F4F532E2E2E2E;
defparam sp_inst_43.INIT_RAM_34 = 256'h2E2E44412E2E2E2E2E2E00002E2E2E2E2E2E2E2E414641422E2E2E2E2E2E0000;
defparam sp_inst_43.INIT_RAM_35 = 256'h6D69657200000A2E7075657420726C63656D20737265697200000A2E2E2E2E2E;
defparam sp_inst_43.INIT_RAM_36 = 256'h1C001C001C001C001C001C001C001C001C001C0000002E2E7572746E72616320;
defparam sp_inst_43.INIT_RAM_37 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_43.INIT_RAM_38 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_43.INIT_RAM_39 = 256'h5F31697069740072646E5F715F30697069741C001C001C001C001C001C001C00;
defparam sp_inst_43.INIT_RAM_3A = 256'h69740072646E5F715F33697069740072646E5F715F32697069740072646E5F71;
defparam sp_inst_43.INIT_RAM_3B = 256'h646E5F715F36697069740072646E5F715F35697069740072646E5F715F346970;
defparam sp_inst_43.INIT_RAM_3C = 256'h5F31697069740072646E5F715F30697069740072646E5F715F37697069740072;
defparam sp_inst_43.INIT_RAM_3D = 256'h69740072646E5F715F33697069740072646E5F715F32697069740072646E5F71;
defparam sp_inst_43.INIT_RAM_3E = 256'h646E5F715F36697069740072646E5F715F35697069740072646E5F715F346970;
defparam sp_inst_43.INIT_RAM_3F = 256'h5F31697069740072646E5F715F30697069740072646E5F715F37697069740072;

SP sp_inst_44 (
    .DO({sp_inst_44_dout_w[15:0],sp_inst_44_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_12}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_44.READ_MODE = 1'b0;
defparam sp_inst_44.WRITE_MODE = 2'b01;
defparam sp_inst_44.BIT_WIDTH = 16;
defparam sp_inst_44.BLK_SEL = 3'b001;
defparam sp_inst_44.RESET_MODE = "SYNC";
defparam sp_inst_44.INIT_RAM_00 = 256'h69740072646E5F715F33697069740072646E5F715F32697069740072646E5F71;
defparam sp_inst_44.INIT_RAM_01 = 256'h646E5F715F36697069740072646E5F715F35697069740072646E5F715F346970;
defparam sp_inst_44.INIT_RAM_02 = 256'h5F31697069740072646E5F715F30697069740072646E5F715F37697069740072;
defparam sp_inst_44.INIT_RAM_03 = 256'h69740072646E5F715F33697069740072646E5F715F32697069740072646E5F71;
defparam sp_inst_44.INIT_RAM_04 = 256'h646E5F715F36697069740072646E5F715F35697069740072646E5F715F346970;
defparam sp_inst_44.INIT_RAM_05 = 256'h8000800080008000800000000072646E5F740072646E5F715F37697069740072;
defparam sp_inst_44.INIT_RAM_06 = 256'h8888007F121200E0888818CC494A0000FF494949FF0000004242105232538000;
defparam sp_inst_44.INIT_RAM_07 = 256'h2909798929490040147F002414240000400000000000000002020202060100E0;
defparam sp_inst_44.INIT_RAM_08 = 256'h3F00304012220088888EC88863AC0000120A7E8213220000810962A232220008;
defparam sp_inst_44.INIT_RAM_09 = 256'hFF0900FF091F0000D20E00E027EC0000080400FF00000040444444FF40400071;
defparam sp_inst_44.INIT_RAM_0A = 256'h43427E42417A000C8414A69504440080100F4F807F01000020BFE200E72C0008;
defparam sp_inst_44.INIT_RAM_0B = 256'hFF0900FF091F0000D20E00E027EC003F48080800107F0080828202005CE40000;
defparam sp_inst_44.INIT_RAM_0C = 256'h462843403F0000209E829EA0CC420080100F4F807F01000020BFE200E72C0008;
defparam sp_inst_44.INIT_RAM_0D = 256'h955515FF207F00405454545400CC00407F5555557F400000D5557D55D5150080;
defparam sp_inst_44.INIT_RAM_0E = 256'h12121212017F00804A524A8610FF0040504F434C1F20000048C8C84ECC420000;
defparam sp_inst_44.INIT_RAM_0F = 256'h100F4F807F01000020BFE200E72C0008FF0900FF091F0000D20E00E027EC0000;
defparam sp_inst_44.INIT_RAM_10 = 256'h100C10102060001010101090909000003F4000002040000888888E8908080080;
defparam sp_inst_44.INIT_RAM_11 = 256'h5F0012FFFF090010941254C8C81F0000955515FF207F00405454545400CC00F8;
defparam sp_inst_44.INIT_RAM_12 = 256'h43427E42417A000C8414A69504440080300C00001020000000001CE200000000;
defparam sp_inst_44.INIT_RAM_13 = 256'hFF0900FF091F0000D20E00E027EC003F48080800107F0080828202005CE40000;
defparam sp_inst_44.INIT_RAM_14 = 256'h21110103214100001010FF101E300080100F4F807F01000020BFE200E72C0008;
defparam sp_inst_44.INIT_RAM_15 = 256'h1816801F001F00080908088888F80080160840800F30001010102040FA020081;
defparam sp_inst_44.INIT_RAM_16 = 256'h4141294500FF00042424242407F80000804030481F10000010101008F80800F8;
defparam sp_inst_44.INIT_RAM_17 = 256'hF84B4A4AFF00006226A2BAA2A223000082427F02021F00002222FE2222FE0080;
defparam sp_inst_44.INIT_RAM_18 = 256'h20200E10408F00005E5252525EC00040447F44401F20000092FEFE00FC840000;
defparam sp_inst_44.INIT_RAM_19 = 256'h40407F40404000004040FF40407C00404241485F1F200000494949FFCC420000;
defparam sp_inst_44.INIT_RAM_1A = 256'h20202424207F00000202121202FE0040454250471F200000222224FCCC420000;
defparam sp_inst_44.INIT_RAM_1B = 256'h427F444F1F20000004FC04FCCC42008018061820010600000808304084440000;
defparam sp_inst_44.INIT_RAM_1C = 256'h213F7F00000000080868182000000078404000002040004048507F4044420040;
defparam sp_inst_44.INIT_RAM_1D = 256'h20202424207F00000202121202FE0040454250471F200000222224FCCC420000;
defparam sp_inst_44.INIT_RAM_1E = 256'h2020007F0F300000080800F0FF10003130084018017E0010523252928C020000;
defparam sp_inst_44.INIT_RAM_1F = 256'h955515FF017E0040545454548C02001012121212100F000424243D6424FC0000;
defparam sp_inst_44.INIT_RAM_20 = 256'h40404040403F0000FE82828282E200000501410D08040020282428105A220000;
defparam sp_inst_44.INIT_RAM_21 = 256'hFC444544FC0000004222FA12828200818989FF811D2100007F4949497F000000;
defparam sp_inst_44.INIT_RAM_22 = 256'h2116214012220000F808F80863AC00004949FF007F82007044443F00FF100001;
defparam sp_inst_44.INIT_RAM_23 = 256'h281084807F810098888E8898FF100000955515FF207F00405454545400CC0080;
defparam sp_inst_44.INIT_RAM_24 = 256'h4949FF007F82007044443F00FF10000202027F82020200002322FC2424240000;
defparam sp_inst_44.INIT_RAM_25 = 256'h300C00001020000000001CE20000004024187F8024220080FE92929292820000;
defparam sp_inst_44.INIT_RAM_26 = 256'h2116214012220000F808F80863AC00004949FF007F82007044443F00FF100080;
defparam sp_inst_44.INIT_RAM_27 = 256'h804030481F10000010101008F80800F81816801F001F00080908088888F80080;
defparam sp_inst_44.INIT_RAM_28 = 256'h160840800F30001010102040FA02008121110103214100001010FF101E300000;
defparam sp_inst_44.INIT_RAM_29 = 256'h2212FF02023E0018EAACAFA8EA08000808FE0808284800009E929292927E0080;
defparam sp_inst_44.INIT_RAM_2A = 256'h4909FF00FF010000203FE200FEA40000955515FF207F00405454545400CC0000;
defparam sp_inst_44.INIT_RAM_2B = 256'h8444070404FF00029292FE9292F20000424242420718002023222424FC000000;
defparam sp_inst_44.INIT_RAM_2C = 256'h0404FF04040F00001010FF1010F000F00E013F603F00001010FF9090CC420004;
defparam sp_inst_44.INIT_RAM_2D = 256'h80403040FF0000808780B040F86000007F82121223420040FC545455FC000000;
defparam sp_inst_44.INIT_RAM_2E = 256'h417F7F403F00000404FCC404CC420040604E4440844800404C43204082820000;
defparam sp_inst_44.INIT_RAM_2F = 256'h000000000000000000000000000000000000000001E8000000001307FFFF0040;
defparam sp_inst_44.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_45 (
    .DO({sp_inst_45_dout_w[15:0],sp_inst_45_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_13}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_45.READ_MODE = 1'b0;
defparam sp_inst_45.WRITE_MODE = 2'b01;
defparam sp_inst_45.BIT_WIDTH = 16;
defparam sp_inst_45.BLK_SEL = 3'b001;
defparam sp_inst_45.RESET_MODE = "SYNC";
defparam sp_inst_45.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_46 (
    .DO({sp_inst_46_dout_w[15:0],sp_inst_46_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_14}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_46.READ_MODE = 1'b0;
defparam sp_inst_46.WRITE_MODE = 2'b01;
defparam sp_inst_46.BIT_WIDTH = 16;
defparam sp_inst_46.BLK_SEL = 3'b001;
defparam sp_inst_46.RESET_MODE = "SYNC";
defparam sp_inst_46.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_47 (
    .DO({sp_inst_47_dout_w[15:0],sp_inst_47_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_15}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_47.READ_MODE = 1'b0;
defparam sp_inst_47.WRITE_MODE = 2'b01;
defparam sp_inst_47.BIT_WIDTH = 16;
defparam sp_inst_47.BLK_SEL = 3'b001;
defparam sp_inst_47.RESET_MODE = "SYNC";
defparam sp_inst_47.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_48 (
    .DO({sp_inst_48_dout_w[15:0],sp_inst_48_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_16}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_48.READ_MODE = 1'b0;
defparam sp_inst_48.WRITE_MODE = 2'b01;
defparam sp_inst_48.BIT_WIDTH = 16;
defparam sp_inst_48.BLK_SEL = 3'b001;
defparam sp_inst_48.RESET_MODE = "SYNC";
defparam sp_inst_48.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_49 (
    .DO({sp_inst_49_dout_w[15:0],sp_inst_49_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_17}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_49.READ_MODE = 1'b0;
defparam sp_inst_49.WRITE_MODE = 2'b01;
defparam sp_inst_49.BIT_WIDTH = 16;
defparam sp_inst_49.BLK_SEL = 3'b001;
defparam sp_inst_49.RESET_MODE = "SYNC";
defparam sp_inst_49.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_50 (
    .DO({sp_inst_50_dout_w[15:0],sp_inst_50_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_18}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_50.READ_MODE = 1'b0;
defparam sp_inst_50.WRITE_MODE = 2'b01;
defparam sp_inst_50.BIT_WIDTH = 16;
defparam sp_inst_50.BLK_SEL = 3'b001;
defparam sp_inst_50.RESET_MODE = "SYNC";
defparam sp_inst_50.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_51 (
    .DO({sp_inst_51_dout_w[15:0],sp_inst_51_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_19}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_51.READ_MODE = 1'b0;
defparam sp_inst_51.WRITE_MODE = 2'b01;
defparam sp_inst_51.BIT_WIDTH = 16;
defparam sp_inst_51.BLK_SEL = 3'b001;
defparam sp_inst_51.RESET_MODE = "SYNC";
defparam sp_inst_51.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_52 (
    .DO({sp_inst_52_dout_w[15:0],sp_inst_52_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_20}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_52.READ_MODE = 1'b0;
defparam sp_inst_52.WRITE_MODE = 2'b01;
defparam sp_inst_52.BIT_WIDTH = 16;
defparam sp_inst_52.BLK_SEL = 3'b001;
defparam sp_inst_52.RESET_MODE = "SYNC";
defparam sp_inst_52.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_53 (
    .DO({sp_inst_53_dout_w[15:0],sp_inst_53_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_21}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_53.READ_MODE = 1'b0;
defparam sp_inst_53.WRITE_MODE = 2'b01;
defparam sp_inst_53.BIT_WIDTH = 16;
defparam sp_inst_53.BLK_SEL = 3'b001;
defparam sp_inst_53.RESET_MODE = "SYNC";
defparam sp_inst_53.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_54 (
    .DO({sp_inst_54_dout_w[15:0],sp_inst_54_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_22}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_54.READ_MODE = 1'b0;
defparam sp_inst_54.WRITE_MODE = 2'b01;
defparam sp_inst_54.BIT_WIDTH = 16;
defparam sp_inst_54.BLK_SEL = 3'b001;
defparam sp_inst_54.RESET_MODE = "SYNC";
defparam sp_inst_54.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_55 (
    .DO({sp_inst_55_dout_w[15:0],sp_inst_55_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_23}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_55.READ_MODE = 1'b0;
defparam sp_inst_55.WRITE_MODE = 2'b01;
defparam sp_inst_55.BIT_WIDTH = 16;
defparam sp_inst_55.BLK_SEL = 3'b001;
defparam sp_inst_55.RESET_MODE = "SYNC";
defparam sp_inst_55.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_56 (
    .DO({sp_inst_56_dout_w[15:0],sp_inst_56_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_24}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_56.READ_MODE = 1'b0;
defparam sp_inst_56.WRITE_MODE = 2'b01;
defparam sp_inst_56.BIT_WIDTH = 16;
defparam sp_inst_56.BLK_SEL = 3'b001;
defparam sp_inst_56.RESET_MODE = "SYNC";
defparam sp_inst_56.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_57 (
    .DO({sp_inst_57_dout_w[15:0],sp_inst_57_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_25}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_57.READ_MODE = 1'b0;
defparam sp_inst_57.WRITE_MODE = 2'b01;
defparam sp_inst_57.BIT_WIDTH = 16;
defparam sp_inst_57.BLK_SEL = 3'b001;
defparam sp_inst_57.RESET_MODE = "SYNC";
defparam sp_inst_57.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_58 (
    .DO({sp_inst_58_dout_w[15:0],sp_inst_58_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_26}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_58.READ_MODE = 1'b0;
defparam sp_inst_58.WRITE_MODE = 2'b01;
defparam sp_inst_58.BIT_WIDTH = 16;
defparam sp_inst_58.BLK_SEL = 3'b001;
defparam sp_inst_58.RESET_MODE = "SYNC";
defparam sp_inst_58.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_59 (
    .DO({sp_inst_59_dout_w[15:0],sp_inst_59_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_27}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_59.READ_MODE = 1'b0;
defparam sp_inst_59.WRITE_MODE = 2'b01;
defparam sp_inst_59.BIT_WIDTH = 16;
defparam sp_inst_59.BLK_SEL = 3'b001;
defparam sp_inst_59.RESET_MODE = "SYNC";
defparam sp_inst_59.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_60 (
    .DO({sp_inst_60_dout_w[15:0],sp_inst_60_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_28}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_60.READ_MODE = 1'b0;
defparam sp_inst_60.WRITE_MODE = 2'b01;
defparam sp_inst_60.BIT_WIDTH = 16;
defparam sp_inst_60.BLK_SEL = 3'b001;
defparam sp_inst_60.RESET_MODE = "SYNC";
defparam sp_inst_60.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_61 (
    .DO({sp_inst_61_dout_w[15:0],sp_inst_61_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_29}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_61.READ_MODE = 1'b0;
defparam sp_inst_61.WRITE_MODE = 2'b01;
defparam sp_inst_61.BIT_WIDTH = 16;
defparam sp_inst_61.BLK_SEL = 3'b001;
defparam sp_inst_61.RESET_MODE = "SYNC";
defparam sp_inst_61.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_62 (
    .DO({sp_inst_62_dout_w[15:0],sp_inst_62_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_30}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_62.READ_MODE = 1'b0;
defparam sp_inst_62.WRITE_MODE = 2'b01;
defparam sp_inst_62.BIT_WIDTH = 16;
defparam sp_inst_62.BLK_SEL = 3'b001;
defparam sp_inst_62.RESET_MODE = "SYNC";
defparam sp_inst_62.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_63 (
    .DO({sp_inst_63_dout_w[15:0],sp_inst_63_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_31}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_63.READ_MODE = 1'b0;
defparam sp_inst_63.WRITE_MODE = 2'b01;
defparam sp_inst_63.BIT_WIDTH = 16;
defparam sp_inst_63.BLK_SEL = 3'b001;
defparam sp_inst_63.RESET_MODE = "SYNC";
defparam sp_inst_63.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
DFFRE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
DFFRE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
DFFRE dff_inst_3 (
  .Q(dff_q_3),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
DFFRE dff_inst_4 (
  .Q(dff_q_4),
  .D(ad[10]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(sp_inst_0_dout[0]),
  .I1(sp_inst_1_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(sp_inst_2_dout[0]),
  .I1(sp_inst_3_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(sp_inst_4_dout[0]),
  .I1(sp_inst_5_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(sp_inst_6_dout[0]),
  .I1(sp_inst_7_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(sp_inst_8_dout[0]),
  .I1(sp_inst_9_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(sp_inst_10_dout[0]),
  .I1(sp_inst_11_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(sp_inst_12_dout[0]),
  .I1(sp_inst_13_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(sp_inst_14_dout[0]),
  .I1(sp_inst_15_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(sp_inst_16_dout[0]),
  .I1(sp_inst_17_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(sp_inst_18_dout[0]),
  .I1(sp_inst_19_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(sp_inst_20_dout[0]),
  .I1(sp_inst_21_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(sp_inst_22_dout[0]),
  .I1(sp_inst_23_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(sp_inst_24_dout[0]),
  .I1(sp_inst_25_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(sp_inst_26_dout[0]),
  .I1(sp_inst_27_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(sp_inst_28_dout[0]),
  .I1(sp_inst_29_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(sp_inst_30_dout[0]),
  .I1(sp_inst_31_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_3)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_3)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_3)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(dff_q_3)
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(dff_q_3)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_3)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_3)
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(dff_q_3)
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(dff_q_2)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(dff_q_2)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(mux_o_20),
  .I1(mux_o_21),
  .S0(dff_q_2)
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(mux_o_22),
  .I1(mux_o_23),
  .S0(dff_q_2)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(mux_o_24),
  .I1(mux_o_25),
  .S0(dff_q_1)
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(mux_o_26),
  .I1(mux_o_27),
  .S0(dff_q_1)
);
MUX2 mux_inst_30 (
  .O(dout[0]),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(dff_q_0)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(sp_inst_0_dout[1]),
  .I1(sp_inst_1_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(sp_inst_2_dout[1]),
  .I1(sp_inst_3_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(sp_inst_4_dout[1]),
  .I1(sp_inst_5_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(sp_inst_6_dout[1]),
  .I1(sp_inst_7_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(sp_inst_8_dout[1]),
  .I1(sp_inst_9_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(sp_inst_10_dout[1]),
  .I1(sp_inst_11_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(sp_inst_12_dout[1]),
  .I1(sp_inst_13_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(sp_inst_14_dout[1]),
  .I1(sp_inst_15_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(sp_inst_16_dout[1]),
  .I1(sp_inst_17_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(sp_inst_18_dout[1]),
  .I1(sp_inst_19_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(sp_inst_20_dout[1]),
  .I1(sp_inst_21_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(sp_inst_22_dout[1]),
  .I1(sp_inst_23_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(sp_inst_24_dout[1]),
  .I1(sp_inst_25_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(sp_inst_26_dout[1]),
  .I1(sp_inst_27_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(sp_inst_28_dout[1]),
  .I1(sp_inst_29_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(sp_inst_30_dout[1]),
  .I1(sp_inst_31_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(mux_o_31),
  .I1(mux_o_32),
  .S0(dff_q_3)
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(mux_o_33),
  .I1(mux_o_34),
  .S0(dff_q_3)
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(mux_o_35),
  .I1(mux_o_36),
  .S0(dff_q_3)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(mux_o_37),
  .I1(mux_o_38),
  .S0(dff_q_3)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(mux_o_39),
  .I1(mux_o_40),
  .S0(dff_q_3)
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(mux_o_41),
  .I1(mux_o_42),
  .S0(dff_q_3)
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_43),
  .I1(mux_o_44),
  .S0(dff_q_3)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(dff_q_3)
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(mux_o_47),
  .I1(mux_o_48),
  .S0(dff_q_2)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(dff_q_2)
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(mux_o_51),
  .I1(mux_o_52),
  .S0(dff_q_2)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(mux_o_53),
  .I1(mux_o_54),
  .S0(dff_q_2)
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(mux_o_55),
  .I1(mux_o_56),
  .S0(dff_q_1)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(mux_o_57),
  .I1(mux_o_58),
  .S0(dff_q_1)
);
MUX2 mux_inst_61 (
  .O(dout[1]),
  .I0(mux_o_59),
  .I1(mux_o_60),
  .S0(dff_q_0)
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(sp_inst_0_dout[2]),
  .I1(sp_inst_1_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(sp_inst_2_dout[2]),
  .I1(sp_inst_3_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(sp_inst_4_dout[2]),
  .I1(sp_inst_5_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(sp_inst_6_dout[2]),
  .I1(sp_inst_7_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(sp_inst_8_dout[2]),
  .I1(sp_inst_9_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(sp_inst_10_dout[2]),
  .I1(sp_inst_11_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(sp_inst_12_dout[2]),
  .I1(sp_inst_13_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(sp_inst_14_dout[2]),
  .I1(sp_inst_15_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(sp_inst_16_dout[2]),
  .I1(sp_inst_17_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(sp_inst_18_dout[2]),
  .I1(sp_inst_19_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(sp_inst_20_dout[2]),
  .I1(sp_inst_21_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(sp_inst_22_dout[2]),
  .I1(sp_inst_23_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(sp_inst_24_dout[2]),
  .I1(sp_inst_25_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(sp_inst_26_dout[2]),
  .I1(sp_inst_27_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(sp_inst_28_dout[2]),
  .I1(sp_inst_29_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(sp_inst_30_dout[2]),
  .I1(sp_inst_31_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(dff_q_3)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(mux_o_64),
  .I1(mux_o_65),
  .S0(dff_q_3)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(dff_q_3)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(mux_o_68),
  .I1(mux_o_69),
  .S0(dff_q_3)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(dff_q_3)
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(dff_q_3)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(mux_o_74),
  .I1(mux_o_75),
  .S0(dff_q_3)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(mux_o_76),
  .I1(mux_o_77),
  .S0(dff_q_3)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(mux_o_78),
  .I1(mux_o_79),
  .S0(dff_q_2)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(mux_o_80),
  .I1(mux_o_81),
  .S0(dff_q_2)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_82),
  .I1(mux_o_83),
  .S0(dff_q_2)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(mux_o_84),
  .I1(mux_o_85),
  .S0(dff_q_2)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(mux_o_86),
  .I1(mux_o_87),
  .S0(dff_q_1)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(mux_o_88),
  .I1(mux_o_89),
  .S0(dff_q_1)
);
MUX2 mux_inst_92 (
  .O(dout[2]),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(dff_q_0)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(sp_inst_0_dout[3]),
  .I1(sp_inst_1_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(sp_inst_2_dout[3]),
  .I1(sp_inst_3_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(sp_inst_4_dout[3]),
  .I1(sp_inst_5_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(sp_inst_6_dout[3]),
  .I1(sp_inst_7_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(sp_inst_8_dout[3]),
  .I1(sp_inst_9_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(sp_inst_10_dout[3]),
  .I1(sp_inst_11_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(sp_inst_12_dout[3]),
  .I1(sp_inst_13_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(sp_inst_14_dout[3]),
  .I1(sp_inst_15_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(sp_inst_16_dout[3]),
  .I1(sp_inst_17_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(sp_inst_18_dout[3]),
  .I1(sp_inst_19_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(sp_inst_20_dout[3]),
  .I1(sp_inst_21_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_104 (
  .O(mux_o_104),
  .I0(sp_inst_22_dout[3]),
  .I1(sp_inst_23_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(sp_inst_24_dout[3]),
  .I1(sp_inst_25_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(sp_inst_26_dout[3]),
  .I1(sp_inst_27_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(sp_inst_28_dout[3]),
  .I1(sp_inst_29_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(sp_inst_30_dout[3]),
  .I1(sp_inst_31_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(mux_o_93),
  .I1(mux_o_94),
  .S0(dff_q_3)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(mux_o_95),
  .I1(mux_o_96),
  .S0(dff_q_3)
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(mux_o_97),
  .I1(mux_o_98),
  .S0(dff_q_3)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(mux_o_99),
  .I1(mux_o_100),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_101),
  .I1(mux_o_102),
  .S0(dff_q_3)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_103),
  .I1(mux_o_104),
  .S0(dff_q_3)
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(dff_q_3)
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(dff_q_3)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(dff_q_2)
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_111),
  .I1(mux_o_112),
  .S0(dff_q_2)
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(mux_o_113),
  .I1(mux_o_114),
  .S0(dff_q_2)
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(mux_o_115),
  .I1(mux_o_116),
  .S0(dff_q_2)
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(mux_o_117),
  .I1(mux_o_118),
  .S0(dff_q_1)
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(mux_o_119),
  .I1(mux_o_120),
  .S0(dff_q_1)
);
MUX2 mux_inst_123 (
  .O(dout[3]),
  .I0(mux_o_121),
  .I1(mux_o_122),
  .S0(dff_q_0)
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(sp_inst_0_dout[4]),
  .I1(sp_inst_1_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_125 (
  .O(mux_o_125),
  .I0(sp_inst_2_dout[4]),
  .I1(sp_inst_3_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(sp_inst_4_dout[4]),
  .I1(sp_inst_5_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(sp_inst_6_dout[4]),
  .I1(sp_inst_7_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(sp_inst_8_dout[4]),
  .I1(sp_inst_9_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(sp_inst_10_dout[4]),
  .I1(sp_inst_11_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(sp_inst_12_dout[4]),
  .I1(sp_inst_13_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(sp_inst_14_dout[4]),
  .I1(sp_inst_15_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(sp_inst_16_dout[4]),
  .I1(sp_inst_17_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(sp_inst_18_dout[4]),
  .I1(sp_inst_19_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(sp_inst_20_dout[4]),
  .I1(sp_inst_21_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(sp_inst_22_dout[4]),
  .I1(sp_inst_23_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(sp_inst_24_dout[4]),
  .I1(sp_inst_25_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(sp_inst_26_dout[4]),
  .I1(sp_inst_27_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(sp_inst_28_dout[4]),
  .I1(sp_inst_29_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(sp_inst_30_dout[4]),
  .I1(sp_inst_31_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(mux_o_124),
  .I1(mux_o_125),
  .S0(dff_q_3)
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(dff_q_3)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(dff_q_3)
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(dff_q_3)
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(mux_o_132),
  .I1(mux_o_133),
  .S0(dff_q_3)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(mux_o_134),
  .I1(mux_o_135),
  .S0(dff_q_3)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(mux_o_136),
  .I1(mux_o_137),
  .S0(dff_q_3)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(mux_o_138),
  .I1(mux_o_139),
  .S0(dff_q_3)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(mux_o_140),
  .I1(mux_o_141),
  .S0(dff_q_2)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(mux_o_142),
  .I1(mux_o_143),
  .S0(dff_q_2)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(mux_o_144),
  .I1(mux_o_145),
  .S0(dff_q_2)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(mux_o_146),
  .I1(mux_o_147),
  .S0(dff_q_2)
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(mux_o_148),
  .I1(mux_o_149),
  .S0(dff_q_1)
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(mux_o_150),
  .I1(mux_o_151),
  .S0(dff_q_1)
);
MUX2 mux_inst_154 (
  .O(dout[4]),
  .I0(mux_o_152),
  .I1(mux_o_153),
  .S0(dff_q_0)
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(sp_inst_0_dout[5]),
  .I1(sp_inst_1_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(sp_inst_2_dout[5]),
  .I1(sp_inst_3_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(sp_inst_4_dout[5]),
  .I1(sp_inst_5_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(sp_inst_6_dout[5]),
  .I1(sp_inst_7_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(sp_inst_8_dout[5]),
  .I1(sp_inst_9_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(sp_inst_10_dout[5]),
  .I1(sp_inst_11_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(sp_inst_12_dout[5]),
  .I1(sp_inst_13_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(sp_inst_14_dout[5]),
  .I1(sp_inst_15_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(sp_inst_16_dout[5]),
  .I1(sp_inst_17_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(sp_inst_18_dout[5]),
  .I1(sp_inst_19_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(sp_inst_20_dout[5]),
  .I1(sp_inst_21_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(sp_inst_22_dout[5]),
  .I1(sp_inst_23_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(sp_inst_24_dout[5]),
  .I1(sp_inst_25_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(sp_inst_26_dout[5]),
  .I1(sp_inst_27_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(sp_inst_28_dout[5]),
  .I1(sp_inst_29_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(sp_inst_30_dout[5]),
  .I1(sp_inst_31_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(mux_o_155),
  .I1(mux_o_156),
  .S0(dff_q_3)
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(mux_o_157),
  .I1(mux_o_158),
  .S0(dff_q_3)
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(mux_o_159),
  .I1(mux_o_160),
  .S0(dff_q_3)
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(mux_o_161),
  .I1(mux_o_162),
  .S0(dff_q_3)
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(mux_o_163),
  .I1(mux_o_164),
  .S0(dff_q_3)
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(dff_q_3)
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(mux_o_167),
  .I1(mux_o_168),
  .S0(dff_q_3)
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(mux_o_169),
  .I1(mux_o_170),
  .S0(dff_q_3)
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(mux_o_171),
  .I1(mux_o_172),
  .S0(dff_q_2)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(mux_o_173),
  .I1(mux_o_174),
  .S0(dff_q_2)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(mux_o_175),
  .I1(mux_o_176),
  .S0(dff_q_2)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(mux_o_177),
  .I1(mux_o_178),
  .S0(dff_q_2)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(mux_o_179),
  .I1(mux_o_180),
  .S0(dff_q_1)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(mux_o_181),
  .I1(mux_o_182),
  .S0(dff_q_1)
);
MUX2 mux_inst_185 (
  .O(dout[5]),
  .I0(mux_o_183),
  .I1(mux_o_184),
  .S0(dff_q_0)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(sp_inst_0_dout[6]),
  .I1(sp_inst_1_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(sp_inst_2_dout[6]),
  .I1(sp_inst_3_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(sp_inst_4_dout[6]),
  .I1(sp_inst_5_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(sp_inst_6_dout[6]),
  .I1(sp_inst_7_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(sp_inst_8_dout[6]),
  .I1(sp_inst_9_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(sp_inst_10_dout[6]),
  .I1(sp_inst_11_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(sp_inst_12_dout[6]),
  .I1(sp_inst_13_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(sp_inst_14_dout[6]),
  .I1(sp_inst_15_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(sp_inst_16_dout[6]),
  .I1(sp_inst_17_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(sp_inst_18_dout[6]),
  .I1(sp_inst_19_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(sp_inst_20_dout[6]),
  .I1(sp_inst_21_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(sp_inst_22_dout[6]),
  .I1(sp_inst_23_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(sp_inst_24_dout[6]),
  .I1(sp_inst_25_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(sp_inst_26_dout[6]),
  .I1(sp_inst_27_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(sp_inst_28_dout[6]),
  .I1(sp_inst_29_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(sp_inst_30_dout[6]),
  .I1(sp_inst_31_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(dff_q_3)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_188),
  .I1(mux_o_189),
  .S0(dff_q_3)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(mux_o_190),
  .I1(mux_o_191),
  .S0(dff_q_3)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_192),
  .I1(mux_o_193),
  .S0(dff_q_3)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_194),
  .I1(mux_o_195),
  .S0(dff_q_3)
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(mux_o_196),
  .I1(mux_o_197),
  .S0(dff_q_3)
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(mux_o_198),
  .I1(mux_o_199),
  .S0(dff_q_3)
);
MUX2 mux_inst_209 (
  .O(mux_o_209),
  .I0(mux_o_200),
  .I1(mux_o_201),
  .S0(dff_q_3)
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(mux_o_202),
  .I1(mux_o_203),
  .S0(dff_q_2)
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(mux_o_204),
  .I1(mux_o_205),
  .S0(dff_q_2)
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(mux_o_206),
  .I1(mux_o_207),
  .S0(dff_q_2)
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(mux_o_208),
  .I1(mux_o_209),
  .S0(dff_q_2)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(mux_o_210),
  .I1(mux_o_211),
  .S0(dff_q_1)
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(mux_o_212),
  .I1(mux_o_213),
  .S0(dff_q_1)
);
MUX2 mux_inst_216 (
  .O(dout[6]),
  .I0(mux_o_214),
  .I1(mux_o_215),
  .S0(dff_q_0)
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(sp_inst_0_dout[7]),
  .I1(sp_inst_1_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(sp_inst_2_dout[7]),
  .I1(sp_inst_3_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(sp_inst_4_dout[7]),
  .I1(sp_inst_5_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(sp_inst_6_dout[7]),
  .I1(sp_inst_7_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(sp_inst_8_dout[7]),
  .I1(sp_inst_9_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(sp_inst_10_dout[7]),
  .I1(sp_inst_11_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(sp_inst_12_dout[7]),
  .I1(sp_inst_13_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(sp_inst_14_dout[7]),
  .I1(sp_inst_15_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(sp_inst_16_dout[7]),
  .I1(sp_inst_17_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(sp_inst_18_dout[7]),
  .I1(sp_inst_19_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(sp_inst_20_dout[7]),
  .I1(sp_inst_21_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(sp_inst_22_dout[7]),
  .I1(sp_inst_23_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(sp_inst_24_dout[7]),
  .I1(sp_inst_25_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(sp_inst_26_dout[7]),
  .I1(sp_inst_27_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(sp_inst_28_dout[7]),
  .I1(sp_inst_29_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(sp_inst_30_dout[7]),
  .I1(sp_inst_31_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_217),
  .I1(mux_o_218),
  .S0(dff_q_3)
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(mux_o_219),
  .I1(mux_o_220),
  .S0(dff_q_3)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_221),
  .I1(mux_o_222),
  .S0(dff_q_3)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_223),
  .I1(mux_o_224),
  .S0(dff_q_3)
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_225),
  .I1(mux_o_226),
  .S0(dff_q_3)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_227),
  .I1(mux_o_228),
  .S0(dff_q_3)
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(mux_o_229),
  .I1(mux_o_230),
  .S0(dff_q_3)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(dff_q_3)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(dff_q_2)
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_2)
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(dff_q_2)
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(mux_o_239),
  .I1(mux_o_240),
  .S0(dff_q_2)
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(mux_o_241),
  .I1(mux_o_242),
  .S0(dff_q_1)
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(mux_o_243),
  .I1(mux_o_244),
  .S0(dff_q_1)
);
MUX2 mux_inst_247 (
  .O(dout[7]),
  .I0(mux_o_245),
  .I1(mux_o_246),
  .S0(dff_q_0)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(sp_inst_0_dout[8]),
  .I1(sp_inst_1_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(sp_inst_2_dout[8]),
  .I1(sp_inst_3_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(sp_inst_4_dout[8]),
  .I1(sp_inst_5_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_251 (
  .O(mux_o_251),
  .I0(sp_inst_6_dout[8]),
  .I1(sp_inst_7_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(sp_inst_8_dout[8]),
  .I1(sp_inst_9_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(sp_inst_10_dout[8]),
  .I1(sp_inst_11_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(sp_inst_12_dout[8]),
  .I1(sp_inst_13_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(sp_inst_14_dout[8]),
  .I1(sp_inst_15_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(sp_inst_16_dout[8]),
  .I1(sp_inst_17_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(sp_inst_18_dout[8]),
  .I1(sp_inst_19_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(sp_inst_20_dout[8]),
  .I1(sp_inst_21_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(sp_inst_22_dout[8]),
  .I1(sp_inst_23_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(sp_inst_24_dout[8]),
  .I1(sp_inst_25_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(sp_inst_26_dout[8]),
  .I1(sp_inst_27_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(sp_inst_28_dout[8]),
  .I1(sp_inst_29_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(sp_inst_30_dout[8]),
  .I1(sp_inst_31_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(mux_o_248),
  .I1(mux_o_249),
  .S0(dff_q_3)
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(mux_o_250),
  .I1(mux_o_251),
  .S0(dff_q_3)
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(mux_o_252),
  .I1(mux_o_253),
  .S0(dff_q_3)
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(mux_o_254),
  .I1(mux_o_255),
  .S0(dff_q_3)
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(mux_o_256),
  .I1(mux_o_257),
  .S0(dff_q_3)
);
MUX2 mux_inst_269 (
  .O(mux_o_269),
  .I0(mux_o_258),
  .I1(mux_o_259),
  .S0(dff_q_3)
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(mux_o_260),
  .I1(mux_o_261),
  .S0(dff_q_3)
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(mux_o_262),
  .I1(mux_o_263),
  .S0(dff_q_3)
);
MUX2 mux_inst_272 (
  .O(mux_o_272),
  .I0(mux_o_264),
  .I1(mux_o_265),
  .S0(dff_q_2)
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(mux_o_266),
  .I1(mux_o_267),
  .S0(dff_q_2)
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(mux_o_268),
  .I1(mux_o_269),
  .S0(dff_q_2)
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(dff_q_2)
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(mux_o_272),
  .I1(mux_o_273),
  .S0(dff_q_1)
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(mux_o_274),
  .I1(mux_o_275),
  .S0(dff_q_1)
);
MUX2 mux_inst_278 (
  .O(dout[8]),
  .I0(mux_o_276),
  .I1(mux_o_277),
  .S0(dff_q_0)
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(sp_inst_0_dout[9]),
  .I1(sp_inst_1_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(sp_inst_2_dout[9]),
  .I1(sp_inst_3_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(sp_inst_4_dout[9]),
  .I1(sp_inst_5_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(sp_inst_6_dout[9]),
  .I1(sp_inst_7_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(sp_inst_8_dout[9]),
  .I1(sp_inst_9_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_284 (
  .O(mux_o_284),
  .I0(sp_inst_10_dout[9]),
  .I1(sp_inst_11_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(sp_inst_12_dout[9]),
  .I1(sp_inst_13_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(sp_inst_14_dout[9]),
  .I1(sp_inst_15_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(sp_inst_16_dout[9]),
  .I1(sp_inst_17_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(sp_inst_18_dout[9]),
  .I1(sp_inst_19_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(sp_inst_20_dout[9]),
  .I1(sp_inst_21_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(sp_inst_22_dout[9]),
  .I1(sp_inst_23_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(sp_inst_24_dout[9]),
  .I1(sp_inst_25_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(sp_inst_26_dout[9]),
  .I1(sp_inst_27_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(sp_inst_28_dout[9]),
  .I1(sp_inst_29_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(sp_inst_30_dout[9]),
  .I1(sp_inst_31_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(mux_o_279),
  .I1(mux_o_280),
  .S0(dff_q_3)
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(mux_o_281),
  .I1(mux_o_282),
  .S0(dff_q_3)
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(mux_o_283),
  .I1(mux_o_284),
  .S0(dff_q_3)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(mux_o_285),
  .I1(mux_o_286),
  .S0(dff_q_3)
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(mux_o_287),
  .I1(mux_o_288),
  .S0(dff_q_3)
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(mux_o_289),
  .I1(mux_o_290),
  .S0(dff_q_3)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(mux_o_291),
  .I1(mux_o_292),
  .S0(dff_q_3)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(mux_o_293),
  .I1(mux_o_294),
  .S0(dff_q_3)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(mux_o_295),
  .I1(mux_o_296),
  .S0(dff_q_2)
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(mux_o_297),
  .I1(mux_o_298),
  .S0(dff_q_2)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(mux_o_299),
  .I1(mux_o_300),
  .S0(dff_q_2)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(mux_o_301),
  .I1(mux_o_302),
  .S0(dff_q_2)
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(mux_o_303),
  .I1(mux_o_304),
  .S0(dff_q_1)
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(mux_o_305),
  .I1(mux_o_306),
  .S0(dff_q_1)
);
MUX2 mux_inst_309 (
  .O(dout[9]),
  .I0(mux_o_307),
  .I1(mux_o_308),
  .S0(dff_q_0)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(sp_inst_0_dout[10]),
  .I1(sp_inst_1_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(sp_inst_2_dout[10]),
  .I1(sp_inst_3_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(sp_inst_4_dout[10]),
  .I1(sp_inst_5_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(sp_inst_6_dout[10]),
  .I1(sp_inst_7_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_314 (
  .O(mux_o_314),
  .I0(sp_inst_8_dout[10]),
  .I1(sp_inst_9_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(sp_inst_10_dout[10]),
  .I1(sp_inst_11_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(sp_inst_12_dout[10]),
  .I1(sp_inst_13_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(sp_inst_14_dout[10]),
  .I1(sp_inst_15_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(sp_inst_16_dout[10]),
  .I1(sp_inst_17_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(sp_inst_18_dout[10]),
  .I1(sp_inst_19_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(sp_inst_20_dout[10]),
  .I1(sp_inst_21_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(sp_inst_22_dout[10]),
  .I1(sp_inst_23_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(sp_inst_24_dout[10]),
  .I1(sp_inst_25_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(sp_inst_26_dout[10]),
  .I1(sp_inst_27_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(sp_inst_28_dout[10]),
  .I1(sp_inst_29_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(sp_inst_30_dout[10]),
  .I1(sp_inst_31_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(dff_q_3)
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(dff_q_3)
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(mux_o_314),
  .I1(mux_o_315),
  .S0(dff_q_3)
);
MUX2 mux_inst_329 (
  .O(mux_o_329),
  .I0(mux_o_316),
  .I1(mux_o_317),
  .S0(dff_q_3)
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(mux_o_318),
  .I1(mux_o_319),
  .S0(dff_q_3)
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(mux_o_320),
  .I1(mux_o_321),
  .S0(dff_q_3)
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(mux_o_322),
  .I1(mux_o_323),
  .S0(dff_q_3)
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(mux_o_324),
  .I1(mux_o_325),
  .S0(dff_q_3)
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(mux_o_326),
  .I1(mux_o_327),
  .S0(dff_q_2)
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(mux_o_328),
  .I1(mux_o_329),
  .S0(dff_q_2)
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(mux_o_330),
  .I1(mux_o_331),
  .S0(dff_q_2)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(mux_o_332),
  .I1(mux_o_333),
  .S0(dff_q_2)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(mux_o_334),
  .I1(mux_o_335),
  .S0(dff_q_1)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(mux_o_336),
  .I1(mux_o_337),
  .S0(dff_q_1)
);
MUX2 mux_inst_340 (
  .O(dout[10]),
  .I0(mux_o_338),
  .I1(mux_o_339),
  .S0(dff_q_0)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(sp_inst_0_dout[11]),
  .I1(sp_inst_1_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(sp_inst_2_dout[11]),
  .I1(sp_inst_3_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(sp_inst_4_dout[11]),
  .I1(sp_inst_5_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(sp_inst_6_dout[11]),
  .I1(sp_inst_7_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(sp_inst_8_dout[11]),
  .I1(sp_inst_9_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(sp_inst_10_dout[11]),
  .I1(sp_inst_11_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(sp_inst_12_dout[11]),
  .I1(sp_inst_13_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(sp_inst_14_dout[11]),
  .I1(sp_inst_15_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_349 (
  .O(mux_o_349),
  .I0(sp_inst_16_dout[11]),
  .I1(sp_inst_17_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(sp_inst_18_dout[11]),
  .I1(sp_inst_19_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(sp_inst_20_dout[11]),
  .I1(sp_inst_21_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(sp_inst_22_dout[11]),
  .I1(sp_inst_23_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(sp_inst_24_dout[11]),
  .I1(sp_inst_25_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(sp_inst_26_dout[11]),
  .I1(sp_inst_27_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(sp_inst_28_dout[11]),
  .I1(sp_inst_29_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_356 (
  .O(mux_o_356),
  .I0(sp_inst_30_dout[11]),
  .I1(sp_inst_31_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_341),
  .I1(mux_o_342),
  .S0(dff_q_3)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_343),
  .I1(mux_o_344),
  .S0(dff_q_3)
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(mux_o_345),
  .I1(mux_o_346),
  .S0(dff_q_3)
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(dff_q_3)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_349),
  .I1(mux_o_350),
  .S0(dff_q_3)
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(mux_o_351),
  .I1(mux_o_352),
  .S0(dff_q_3)
);
MUX2 mux_inst_363 (
  .O(mux_o_363),
  .I0(mux_o_353),
  .I1(mux_o_354),
  .S0(dff_q_3)
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(mux_o_355),
  .I1(mux_o_356),
  .S0(dff_q_3)
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(dff_q_2)
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(mux_o_359),
  .I1(mux_o_360),
  .S0(dff_q_2)
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(mux_o_361),
  .I1(mux_o_362),
  .S0(dff_q_2)
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(mux_o_363),
  .I1(mux_o_364),
  .S0(dff_q_2)
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(mux_o_365),
  .I1(mux_o_366),
  .S0(dff_q_1)
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(mux_o_367),
  .I1(mux_o_368),
  .S0(dff_q_1)
);
MUX2 mux_inst_371 (
  .O(dout[11]),
  .I0(mux_o_369),
  .I1(mux_o_370),
  .S0(dff_q_0)
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(sp_inst_0_dout[12]),
  .I1(sp_inst_1_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(sp_inst_2_dout[12]),
  .I1(sp_inst_3_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_374 (
  .O(mux_o_374),
  .I0(sp_inst_4_dout[12]),
  .I1(sp_inst_5_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(sp_inst_6_dout[12]),
  .I1(sp_inst_7_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(sp_inst_8_dout[12]),
  .I1(sp_inst_9_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_377 (
  .O(mux_o_377),
  .I0(sp_inst_10_dout[12]),
  .I1(sp_inst_11_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_378 (
  .O(mux_o_378),
  .I0(sp_inst_12_dout[12]),
  .I1(sp_inst_13_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_379 (
  .O(mux_o_379),
  .I0(sp_inst_14_dout[12]),
  .I1(sp_inst_15_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_380 (
  .O(mux_o_380),
  .I0(sp_inst_16_dout[12]),
  .I1(sp_inst_17_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_381 (
  .O(mux_o_381),
  .I0(sp_inst_18_dout[12]),
  .I1(sp_inst_19_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_382 (
  .O(mux_o_382),
  .I0(sp_inst_20_dout[12]),
  .I1(sp_inst_21_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_383 (
  .O(mux_o_383),
  .I0(sp_inst_22_dout[12]),
  .I1(sp_inst_23_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_384 (
  .O(mux_o_384),
  .I0(sp_inst_24_dout[12]),
  .I1(sp_inst_25_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(sp_inst_26_dout[12]),
  .I1(sp_inst_27_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_386 (
  .O(mux_o_386),
  .I0(sp_inst_28_dout[12]),
  .I1(sp_inst_29_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_387 (
  .O(mux_o_387),
  .I0(sp_inst_30_dout[12]),
  .I1(sp_inst_31_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(mux_o_372),
  .I1(mux_o_373),
  .S0(dff_q_3)
);
MUX2 mux_inst_389 (
  .O(mux_o_389),
  .I0(mux_o_374),
  .I1(mux_o_375),
  .S0(dff_q_3)
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(mux_o_376),
  .I1(mux_o_377),
  .S0(dff_q_3)
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(mux_o_378),
  .I1(mux_o_379),
  .S0(dff_q_3)
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(mux_o_380),
  .I1(mux_o_381),
  .S0(dff_q_3)
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(mux_o_382),
  .I1(mux_o_383),
  .S0(dff_q_3)
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(mux_o_384),
  .I1(mux_o_385),
  .S0(dff_q_3)
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(mux_o_386),
  .I1(mux_o_387),
  .S0(dff_q_3)
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(mux_o_388),
  .I1(mux_o_389),
  .S0(dff_q_2)
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(mux_o_390),
  .I1(mux_o_391),
  .S0(dff_q_2)
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(mux_o_392),
  .I1(mux_o_393),
  .S0(dff_q_2)
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(mux_o_394),
  .I1(mux_o_395),
  .S0(dff_q_2)
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(mux_o_396),
  .I1(mux_o_397),
  .S0(dff_q_1)
);
MUX2 mux_inst_401 (
  .O(mux_o_401),
  .I0(mux_o_398),
  .I1(mux_o_399),
  .S0(dff_q_1)
);
MUX2 mux_inst_402 (
  .O(dout[12]),
  .I0(mux_o_400),
  .I1(mux_o_401),
  .S0(dff_q_0)
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(sp_inst_0_dout[13]),
  .I1(sp_inst_1_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_404 (
  .O(mux_o_404),
  .I0(sp_inst_2_dout[13]),
  .I1(sp_inst_3_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(sp_inst_4_dout[13]),
  .I1(sp_inst_5_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(sp_inst_6_dout[13]),
  .I1(sp_inst_7_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(sp_inst_8_dout[13]),
  .I1(sp_inst_9_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_408 (
  .O(mux_o_408),
  .I0(sp_inst_10_dout[13]),
  .I1(sp_inst_11_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(sp_inst_12_dout[13]),
  .I1(sp_inst_13_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(sp_inst_14_dout[13]),
  .I1(sp_inst_15_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(sp_inst_16_dout[13]),
  .I1(sp_inst_17_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_412 (
  .O(mux_o_412),
  .I0(sp_inst_18_dout[13]),
  .I1(sp_inst_19_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(sp_inst_20_dout[13]),
  .I1(sp_inst_21_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(sp_inst_22_dout[13]),
  .I1(sp_inst_23_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_415 (
  .O(mux_o_415),
  .I0(sp_inst_24_dout[13]),
  .I1(sp_inst_25_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_416 (
  .O(mux_o_416),
  .I0(sp_inst_26_dout[13]),
  .I1(sp_inst_27_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_417 (
  .O(mux_o_417),
  .I0(sp_inst_28_dout[13]),
  .I1(sp_inst_29_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_418 (
  .O(mux_o_418),
  .I0(sp_inst_30_dout[13]),
  .I1(sp_inst_31_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_419 (
  .O(mux_o_419),
  .I0(mux_o_403),
  .I1(mux_o_404),
  .S0(dff_q_3)
);
MUX2 mux_inst_420 (
  .O(mux_o_420),
  .I0(mux_o_405),
  .I1(mux_o_406),
  .S0(dff_q_3)
);
MUX2 mux_inst_421 (
  .O(mux_o_421),
  .I0(mux_o_407),
  .I1(mux_o_408),
  .S0(dff_q_3)
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(mux_o_409),
  .I1(mux_o_410),
  .S0(dff_q_3)
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(mux_o_411),
  .I1(mux_o_412),
  .S0(dff_q_3)
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(mux_o_413),
  .I1(mux_o_414),
  .S0(dff_q_3)
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(mux_o_415),
  .I1(mux_o_416),
  .S0(dff_q_3)
);
MUX2 mux_inst_426 (
  .O(mux_o_426),
  .I0(mux_o_417),
  .I1(mux_o_418),
  .S0(dff_q_3)
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(mux_o_419),
  .I1(mux_o_420),
  .S0(dff_q_2)
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(mux_o_421),
  .I1(mux_o_422),
  .S0(dff_q_2)
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(mux_o_423),
  .I1(mux_o_424),
  .S0(dff_q_2)
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(mux_o_425),
  .I1(mux_o_426),
  .S0(dff_q_2)
);
MUX2 mux_inst_431 (
  .O(mux_o_431),
  .I0(mux_o_427),
  .I1(mux_o_428),
  .S0(dff_q_1)
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(mux_o_429),
  .I1(mux_o_430),
  .S0(dff_q_1)
);
MUX2 mux_inst_433 (
  .O(dout[13]),
  .I0(mux_o_431),
  .I1(mux_o_432),
  .S0(dff_q_0)
);
MUX2 mux_inst_434 (
  .O(mux_o_434),
  .I0(sp_inst_0_dout[14]),
  .I1(sp_inst_1_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(sp_inst_2_dout[14]),
  .I1(sp_inst_3_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(sp_inst_4_dout[14]),
  .I1(sp_inst_5_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(sp_inst_6_dout[14]),
  .I1(sp_inst_7_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(sp_inst_8_dout[14]),
  .I1(sp_inst_9_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(sp_inst_10_dout[14]),
  .I1(sp_inst_11_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_440 (
  .O(mux_o_440),
  .I0(sp_inst_12_dout[14]),
  .I1(sp_inst_13_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(sp_inst_14_dout[14]),
  .I1(sp_inst_15_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(sp_inst_16_dout[14]),
  .I1(sp_inst_17_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(sp_inst_18_dout[14]),
  .I1(sp_inst_19_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(sp_inst_20_dout[14]),
  .I1(sp_inst_21_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(sp_inst_22_dout[14]),
  .I1(sp_inst_23_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(sp_inst_24_dout[14]),
  .I1(sp_inst_25_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(sp_inst_26_dout[14]),
  .I1(sp_inst_27_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(sp_inst_28_dout[14]),
  .I1(sp_inst_29_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_449 (
  .O(mux_o_449),
  .I0(sp_inst_30_dout[14]),
  .I1(sp_inst_31_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(mux_o_434),
  .I1(mux_o_435),
  .S0(dff_q_3)
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(mux_o_436),
  .I1(mux_o_437),
  .S0(dff_q_3)
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(mux_o_438),
  .I1(mux_o_439),
  .S0(dff_q_3)
);
MUX2 mux_inst_453 (
  .O(mux_o_453),
  .I0(mux_o_440),
  .I1(mux_o_441),
  .S0(dff_q_3)
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(mux_o_442),
  .I1(mux_o_443),
  .S0(dff_q_3)
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(mux_o_444),
  .I1(mux_o_445),
  .S0(dff_q_3)
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(mux_o_446),
  .I1(mux_o_447),
  .S0(dff_q_3)
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(mux_o_448),
  .I1(mux_o_449),
  .S0(dff_q_3)
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(mux_o_450),
  .I1(mux_o_451),
  .S0(dff_q_2)
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(mux_o_452),
  .I1(mux_o_453),
  .S0(dff_q_2)
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(mux_o_454),
  .I1(mux_o_455),
  .S0(dff_q_2)
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(mux_o_456),
  .I1(mux_o_457),
  .S0(dff_q_2)
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(mux_o_458),
  .I1(mux_o_459),
  .S0(dff_q_1)
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(mux_o_460),
  .I1(mux_o_461),
  .S0(dff_q_1)
);
MUX2 mux_inst_464 (
  .O(dout[14]),
  .I0(mux_o_462),
  .I1(mux_o_463),
  .S0(dff_q_0)
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(sp_inst_0_dout[15]),
  .I1(sp_inst_1_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(sp_inst_2_dout[15]),
  .I1(sp_inst_3_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_467 (
  .O(mux_o_467),
  .I0(sp_inst_4_dout[15]),
  .I1(sp_inst_5_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_468 (
  .O(mux_o_468),
  .I0(sp_inst_6_dout[15]),
  .I1(sp_inst_7_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_469 (
  .O(mux_o_469),
  .I0(sp_inst_8_dout[15]),
  .I1(sp_inst_9_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_470 (
  .O(mux_o_470),
  .I0(sp_inst_10_dout[15]),
  .I1(sp_inst_11_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_471 (
  .O(mux_o_471),
  .I0(sp_inst_12_dout[15]),
  .I1(sp_inst_13_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(sp_inst_14_dout[15]),
  .I1(sp_inst_15_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_473 (
  .O(mux_o_473),
  .I0(sp_inst_16_dout[15]),
  .I1(sp_inst_17_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_474 (
  .O(mux_o_474),
  .I0(sp_inst_18_dout[15]),
  .I1(sp_inst_19_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_475 (
  .O(mux_o_475),
  .I0(sp_inst_20_dout[15]),
  .I1(sp_inst_21_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_476 (
  .O(mux_o_476),
  .I0(sp_inst_22_dout[15]),
  .I1(sp_inst_23_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_477 (
  .O(mux_o_477),
  .I0(sp_inst_24_dout[15]),
  .I1(sp_inst_25_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_478 (
  .O(mux_o_478),
  .I0(sp_inst_26_dout[15]),
  .I1(sp_inst_27_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_479 (
  .O(mux_o_479),
  .I0(sp_inst_28_dout[15]),
  .I1(sp_inst_29_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_480 (
  .O(mux_o_480),
  .I0(sp_inst_30_dout[15]),
  .I1(sp_inst_31_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_481 (
  .O(mux_o_481),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(dff_q_3)
);
MUX2 mux_inst_482 (
  .O(mux_o_482),
  .I0(mux_o_467),
  .I1(mux_o_468),
  .S0(dff_q_3)
);
MUX2 mux_inst_483 (
  .O(mux_o_483),
  .I0(mux_o_469),
  .I1(mux_o_470),
  .S0(dff_q_3)
);
MUX2 mux_inst_484 (
  .O(mux_o_484),
  .I0(mux_o_471),
  .I1(mux_o_472),
  .S0(dff_q_3)
);
MUX2 mux_inst_485 (
  .O(mux_o_485),
  .I0(mux_o_473),
  .I1(mux_o_474),
  .S0(dff_q_3)
);
MUX2 mux_inst_486 (
  .O(mux_o_486),
  .I0(mux_o_475),
  .I1(mux_o_476),
  .S0(dff_q_3)
);
MUX2 mux_inst_487 (
  .O(mux_o_487),
  .I0(mux_o_477),
  .I1(mux_o_478),
  .S0(dff_q_3)
);
MUX2 mux_inst_488 (
  .O(mux_o_488),
  .I0(mux_o_479),
  .I1(mux_o_480),
  .S0(dff_q_3)
);
MUX2 mux_inst_489 (
  .O(mux_o_489),
  .I0(mux_o_481),
  .I1(mux_o_482),
  .S0(dff_q_2)
);
MUX2 mux_inst_490 (
  .O(mux_o_490),
  .I0(mux_o_483),
  .I1(mux_o_484),
  .S0(dff_q_2)
);
MUX2 mux_inst_491 (
  .O(mux_o_491),
  .I0(mux_o_485),
  .I1(mux_o_486),
  .S0(dff_q_2)
);
MUX2 mux_inst_492 (
  .O(mux_o_492),
  .I0(mux_o_487),
  .I1(mux_o_488),
  .S0(dff_q_2)
);
MUX2 mux_inst_493 (
  .O(mux_o_493),
  .I0(mux_o_489),
  .I1(mux_o_490),
  .S0(dff_q_1)
);
MUX2 mux_inst_494 (
  .O(mux_o_494),
  .I0(mux_o_491),
  .I1(mux_o_492),
  .S0(dff_q_1)
);
MUX2 mux_inst_495 (
  .O(dout[15]),
  .I0(mux_o_493),
  .I1(mux_o_494),
  .S0(dff_q_0)
);
MUX2 mux_inst_496 (
  .O(mux_o_496),
  .I0(sp_inst_32_dout[16]),
  .I1(sp_inst_33_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_497 (
  .O(mux_o_497),
  .I0(sp_inst_34_dout[16]),
  .I1(sp_inst_35_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_498 (
  .O(mux_o_498),
  .I0(sp_inst_36_dout[16]),
  .I1(sp_inst_37_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_499 (
  .O(mux_o_499),
  .I0(sp_inst_38_dout[16]),
  .I1(sp_inst_39_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_500 (
  .O(mux_o_500),
  .I0(sp_inst_40_dout[16]),
  .I1(sp_inst_41_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_501 (
  .O(mux_o_501),
  .I0(sp_inst_42_dout[16]),
  .I1(sp_inst_43_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_502 (
  .O(mux_o_502),
  .I0(sp_inst_44_dout[16]),
  .I1(sp_inst_45_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_503 (
  .O(mux_o_503),
  .I0(sp_inst_46_dout[16]),
  .I1(sp_inst_47_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_504 (
  .O(mux_o_504),
  .I0(sp_inst_48_dout[16]),
  .I1(sp_inst_49_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_505 (
  .O(mux_o_505),
  .I0(sp_inst_50_dout[16]),
  .I1(sp_inst_51_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_506 (
  .O(mux_o_506),
  .I0(sp_inst_52_dout[16]),
  .I1(sp_inst_53_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_507 (
  .O(mux_o_507),
  .I0(sp_inst_54_dout[16]),
  .I1(sp_inst_55_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_508 (
  .O(mux_o_508),
  .I0(sp_inst_56_dout[16]),
  .I1(sp_inst_57_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_509 (
  .O(mux_o_509),
  .I0(sp_inst_58_dout[16]),
  .I1(sp_inst_59_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_510 (
  .O(mux_o_510),
  .I0(sp_inst_60_dout[16]),
  .I1(sp_inst_61_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_511 (
  .O(mux_o_511),
  .I0(sp_inst_62_dout[16]),
  .I1(sp_inst_63_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_512 (
  .O(mux_o_512),
  .I0(mux_o_496),
  .I1(mux_o_497),
  .S0(dff_q_3)
);
MUX2 mux_inst_513 (
  .O(mux_o_513),
  .I0(mux_o_498),
  .I1(mux_o_499),
  .S0(dff_q_3)
);
MUX2 mux_inst_514 (
  .O(mux_o_514),
  .I0(mux_o_500),
  .I1(mux_o_501),
  .S0(dff_q_3)
);
MUX2 mux_inst_515 (
  .O(mux_o_515),
  .I0(mux_o_502),
  .I1(mux_o_503),
  .S0(dff_q_3)
);
MUX2 mux_inst_516 (
  .O(mux_o_516),
  .I0(mux_o_504),
  .I1(mux_o_505),
  .S0(dff_q_3)
);
MUX2 mux_inst_517 (
  .O(mux_o_517),
  .I0(mux_o_506),
  .I1(mux_o_507),
  .S0(dff_q_3)
);
MUX2 mux_inst_518 (
  .O(mux_o_518),
  .I0(mux_o_508),
  .I1(mux_o_509),
  .S0(dff_q_3)
);
MUX2 mux_inst_519 (
  .O(mux_o_519),
  .I0(mux_o_510),
  .I1(mux_o_511),
  .S0(dff_q_3)
);
MUX2 mux_inst_520 (
  .O(mux_o_520),
  .I0(mux_o_512),
  .I1(mux_o_513),
  .S0(dff_q_2)
);
MUX2 mux_inst_521 (
  .O(mux_o_521),
  .I0(mux_o_514),
  .I1(mux_o_515),
  .S0(dff_q_2)
);
MUX2 mux_inst_522 (
  .O(mux_o_522),
  .I0(mux_o_516),
  .I1(mux_o_517),
  .S0(dff_q_2)
);
MUX2 mux_inst_523 (
  .O(mux_o_523),
  .I0(mux_o_518),
  .I1(mux_o_519),
  .S0(dff_q_2)
);
MUX2 mux_inst_524 (
  .O(mux_o_524),
  .I0(mux_o_520),
  .I1(mux_o_521),
  .S0(dff_q_1)
);
MUX2 mux_inst_525 (
  .O(mux_o_525),
  .I0(mux_o_522),
  .I1(mux_o_523),
  .S0(dff_q_1)
);
MUX2 mux_inst_526 (
  .O(dout[16]),
  .I0(mux_o_524),
  .I1(mux_o_525),
  .S0(dff_q_0)
);
MUX2 mux_inst_527 (
  .O(mux_o_527),
  .I0(sp_inst_32_dout[17]),
  .I1(sp_inst_33_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_528 (
  .O(mux_o_528),
  .I0(sp_inst_34_dout[17]),
  .I1(sp_inst_35_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_529 (
  .O(mux_o_529),
  .I0(sp_inst_36_dout[17]),
  .I1(sp_inst_37_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_530 (
  .O(mux_o_530),
  .I0(sp_inst_38_dout[17]),
  .I1(sp_inst_39_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_531 (
  .O(mux_o_531),
  .I0(sp_inst_40_dout[17]),
  .I1(sp_inst_41_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_532 (
  .O(mux_o_532),
  .I0(sp_inst_42_dout[17]),
  .I1(sp_inst_43_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_533 (
  .O(mux_o_533),
  .I0(sp_inst_44_dout[17]),
  .I1(sp_inst_45_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_534 (
  .O(mux_o_534),
  .I0(sp_inst_46_dout[17]),
  .I1(sp_inst_47_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_535 (
  .O(mux_o_535),
  .I0(sp_inst_48_dout[17]),
  .I1(sp_inst_49_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_536 (
  .O(mux_o_536),
  .I0(sp_inst_50_dout[17]),
  .I1(sp_inst_51_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_537 (
  .O(mux_o_537),
  .I0(sp_inst_52_dout[17]),
  .I1(sp_inst_53_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_538 (
  .O(mux_o_538),
  .I0(sp_inst_54_dout[17]),
  .I1(sp_inst_55_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_539 (
  .O(mux_o_539),
  .I0(sp_inst_56_dout[17]),
  .I1(sp_inst_57_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_540 (
  .O(mux_o_540),
  .I0(sp_inst_58_dout[17]),
  .I1(sp_inst_59_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_541 (
  .O(mux_o_541),
  .I0(sp_inst_60_dout[17]),
  .I1(sp_inst_61_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_542 (
  .O(mux_o_542),
  .I0(sp_inst_62_dout[17]),
  .I1(sp_inst_63_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_543 (
  .O(mux_o_543),
  .I0(mux_o_527),
  .I1(mux_o_528),
  .S0(dff_q_3)
);
MUX2 mux_inst_544 (
  .O(mux_o_544),
  .I0(mux_o_529),
  .I1(mux_o_530),
  .S0(dff_q_3)
);
MUX2 mux_inst_545 (
  .O(mux_o_545),
  .I0(mux_o_531),
  .I1(mux_o_532),
  .S0(dff_q_3)
);
MUX2 mux_inst_546 (
  .O(mux_o_546),
  .I0(mux_o_533),
  .I1(mux_o_534),
  .S0(dff_q_3)
);
MUX2 mux_inst_547 (
  .O(mux_o_547),
  .I0(mux_o_535),
  .I1(mux_o_536),
  .S0(dff_q_3)
);
MUX2 mux_inst_548 (
  .O(mux_o_548),
  .I0(mux_o_537),
  .I1(mux_o_538),
  .S0(dff_q_3)
);
MUX2 mux_inst_549 (
  .O(mux_o_549),
  .I0(mux_o_539),
  .I1(mux_o_540),
  .S0(dff_q_3)
);
MUX2 mux_inst_550 (
  .O(mux_o_550),
  .I0(mux_o_541),
  .I1(mux_o_542),
  .S0(dff_q_3)
);
MUX2 mux_inst_551 (
  .O(mux_o_551),
  .I0(mux_o_543),
  .I1(mux_o_544),
  .S0(dff_q_2)
);
MUX2 mux_inst_552 (
  .O(mux_o_552),
  .I0(mux_o_545),
  .I1(mux_o_546),
  .S0(dff_q_2)
);
MUX2 mux_inst_553 (
  .O(mux_o_553),
  .I0(mux_o_547),
  .I1(mux_o_548),
  .S0(dff_q_2)
);
MUX2 mux_inst_554 (
  .O(mux_o_554),
  .I0(mux_o_549),
  .I1(mux_o_550),
  .S0(dff_q_2)
);
MUX2 mux_inst_555 (
  .O(mux_o_555),
  .I0(mux_o_551),
  .I1(mux_o_552),
  .S0(dff_q_1)
);
MUX2 mux_inst_556 (
  .O(mux_o_556),
  .I0(mux_o_553),
  .I1(mux_o_554),
  .S0(dff_q_1)
);
MUX2 mux_inst_557 (
  .O(dout[17]),
  .I0(mux_o_555),
  .I1(mux_o_556),
  .S0(dff_q_0)
);
MUX2 mux_inst_558 (
  .O(mux_o_558),
  .I0(sp_inst_32_dout[18]),
  .I1(sp_inst_33_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_559 (
  .O(mux_o_559),
  .I0(sp_inst_34_dout[18]),
  .I1(sp_inst_35_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_560 (
  .O(mux_o_560),
  .I0(sp_inst_36_dout[18]),
  .I1(sp_inst_37_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_561 (
  .O(mux_o_561),
  .I0(sp_inst_38_dout[18]),
  .I1(sp_inst_39_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_562 (
  .O(mux_o_562),
  .I0(sp_inst_40_dout[18]),
  .I1(sp_inst_41_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_563 (
  .O(mux_o_563),
  .I0(sp_inst_42_dout[18]),
  .I1(sp_inst_43_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_564 (
  .O(mux_o_564),
  .I0(sp_inst_44_dout[18]),
  .I1(sp_inst_45_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_565 (
  .O(mux_o_565),
  .I0(sp_inst_46_dout[18]),
  .I1(sp_inst_47_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_566 (
  .O(mux_o_566),
  .I0(sp_inst_48_dout[18]),
  .I1(sp_inst_49_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_567 (
  .O(mux_o_567),
  .I0(sp_inst_50_dout[18]),
  .I1(sp_inst_51_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_568 (
  .O(mux_o_568),
  .I0(sp_inst_52_dout[18]),
  .I1(sp_inst_53_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_569 (
  .O(mux_o_569),
  .I0(sp_inst_54_dout[18]),
  .I1(sp_inst_55_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_570 (
  .O(mux_o_570),
  .I0(sp_inst_56_dout[18]),
  .I1(sp_inst_57_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_571 (
  .O(mux_o_571),
  .I0(sp_inst_58_dout[18]),
  .I1(sp_inst_59_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_572 (
  .O(mux_o_572),
  .I0(sp_inst_60_dout[18]),
  .I1(sp_inst_61_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_573 (
  .O(mux_o_573),
  .I0(sp_inst_62_dout[18]),
  .I1(sp_inst_63_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_574 (
  .O(mux_o_574),
  .I0(mux_o_558),
  .I1(mux_o_559),
  .S0(dff_q_3)
);
MUX2 mux_inst_575 (
  .O(mux_o_575),
  .I0(mux_o_560),
  .I1(mux_o_561),
  .S0(dff_q_3)
);
MUX2 mux_inst_576 (
  .O(mux_o_576),
  .I0(mux_o_562),
  .I1(mux_o_563),
  .S0(dff_q_3)
);
MUX2 mux_inst_577 (
  .O(mux_o_577),
  .I0(mux_o_564),
  .I1(mux_o_565),
  .S0(dff_q_3)
);
MUX2 mux_inst_578 (
  .O(mux_o_578),
  .I0(mux_o_566),
  .I1(mux_o_567),
  .S0(dff_q_3)
);
MUX2 mux_inst_579 (
  .O(mux_o_579),
  .I0(mux_o_568),
  .I1(mux_o_569),
  .S0(dff_q_3)
);
MUX2 mux_inst_580 (
  .O(mux_o_580),
  .I0(mux_o_570),
  .I1(mux_o_571),
  .S0(dff_q_3)
);
MUX2 mux_inst_581 (
  .O(mux_o_581),
  .I0(mux_o_572),
  .I1(mux_o_573),
  .S0(dff_q_3)
);
MUX2 mux_inst_582 (
  .O(mux_o_582),
  .I0(mux_o_574),
  .I1(mux_o_575),
  .S0(dff_q_2)
);
MUX2 mux_inst_583 (
  .O(mux_o_583),
  .I0(mux_o_576),
  .I1(mux_o_577),
  .S0(dff_q_2)
);
MUX2 mux_inst_584 (
  .O(mux_o_584),
  .I0(mux_o_578),
  .I1(mux_o_579),
  .S0(dff_q_2)
);
MUX2 mux_inst_585 (
  .O(mux_o_585),
  .I0(mux_o_580),
  .I1(mux_o_581),
  .S0(dff_q_2)
);
MUX2 mux_inst_586 (
  .O(mux_o_586),
  .I0(mux_o_582),
  .I1(mux_o_583),
  .S0(dff_q_1)
);
MUX2 mux_inst_587 (
  .O(mux_o_587),
  .I0(mux_o_584),
  .I1(mux_o_585),
  .S0(dff_q_1)
);
MUX2 mux_inst_588 (
  .O(dout[18]),
  .I0(mux_o_586),
  .I1(mux_o_587),
  .S0(dff_q_0)
);
MUX2 mux_inst_589 (
  .O(mux_o_589),
  .I0(sp_inst_32_dout[19]),
  .I1(sp_inst_33_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_590 (
  .O(mux_o_590),
  .I0(sp_inst_34_dout[19]),
  .I1(sp_inst_35_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_591 (
  .O(mux_o_591),
  .I0(sp_inst_36_dout[19]),
  .I1(sp_inst_37_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_592 (
  .O(mux_o_592),
  .I0(sp_inst_38_dout[19]),
  .I1(sp_inst_39_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_593 (
  .O(mux_o_593),
  .I0(sp_inst_40_dout[19]),
  .I1(sp_inst_41_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_594 (
  .O(mux_o_594),
  .I0(sp_inst_42_dout[19]),
  .I1(sp_inst_43_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_595 (
  .O(mux_o_595),
  .I0(sp_inst_44_dout[19]),
  .I1(sp_inst_45_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_596 (
  .O(mux_o_596),
  .I0(sp_inst_46_dout[19]),
  .I1(sp_inst_47_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_597 (
  .O(mux_o_597),
  .I0(sp_inst_48_dout[19]),
  .I1(sp_inst_49_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_598 (
  .O(mux_o_598),
  .I0(sp_inst_50_dout[19]),
  .I1(sp_inst_51_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_599 (
  .O(mux_o_599),
  .I0(sp_inst_52_dout[19]),
  .I1(sp_inst_53_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_600 (
  .O(mux_o_600),
  .I0(sp_inst_54_dout[19]),
  .I1(sp_inst_55_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_601 (
  .O(mux_o_601),
  .I0(sp_inst_56_dout[19]),
  .I1(sp_inst_57_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_602 (
  .O(mux_o_602),
  .I0(sp_inst_58_dout[19]),
  .I1(sp_inst_59_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_603 (
  .O(mux_o_603),
  .I0(sp_inst_60_dout[19]),
  .I1(sp_inst_61_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_604 (
  .O(mux_o_604),
  .I0(sp_inst_62_dout[19]),
  .I1(sp_inst_63_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_605 (
  .O(mux_o_605),
  .I0(mux_o_589),
  .I1(mux_o_590),
  .S0(dff_q_3)
);
MUX2 mux_inst_606 (
  .O(mux_o_606),
  .I0(mux_o_591),
  .I1(mux_o_592),
  .S0(dff_q_3)
);
MUX2 mux_inst_607 (
  .O(mux_o_607),
  .I0(mux_o_593),
  .I1(mux_o_594),
  .S0(dff_q_3)
);
MUX2 mux_inst_608 (
  .O(mux_o_608),
  .I0(mux_o_595),
  .I1(mux_o_596),
  .S0(dff_q_3)
);
MUX2 mux_inst_609 (
  .O(mux_o_609),
  .I0(mux_o_597),
  .I1(mux_o_598),
  .S0(dff_q_3)
);
MUX2 mux_inst_610 (
  .O(mux_o_610),
  .I0(mux_o_599),
  .I1(mux_o_600),
  .S0(dff_q_3)
);
MUX2 mux_inst_611 (
  .O(mux_o_611),
  .I0(mux_o_601),
  .I1(mux_o_602),
  .S0(dff_q_3)
);
MUX2 mux_inst_612 (
  .O(mux_o_612),
  .I0(mux_o_603),
  .I1(mux_o_604),
  .S0(dff_q_3)
);
MUX2 mux_inst_613 (
  .O(mux_o_613),
  .I0(mux_o_605),
  .I1(mux_o_606),
  .S0(dff_q_2)
);
MUX2 mux_inst_614 (
  .O(mux_o_614),
  .I0(mux_o_607),
  .I1(mux_o_608),
  .S0(dff_q_2)
);
MUX2 mux_inst_615 (
  .O(mux_o_615),
  .I0(mux_o_609),
  .I1(mux_o_610),
  .S0(dff_q_2)
);
MUX2 mux_inst_616 (
  .O(mux_o_616),
  .I0(mux_o_611),
  .I1(mux_o_612),
  .S0(dff_q_2)
);
MUX2 mux_inst_617 (
  .O(mux_o_617),
  .I0(mux_o_613),
  .I1(mux_o_614),
  .S0(dff_q_1)
);
MUX2 mux_inst_618 (
  .O(mux_o_618),
  .I0(mux_o_615),
  .I1(mux_o_616),
  .S0(dff_q_1)
);
MUX2 mux_inst_619 (
  .O(dout[19]),
  .I0(mux_o_617),
  .I1(mux_o_618),
  .S0(dff_q_0)
);
MUX2 mux_inst_620 (
  .O(mux_o_620),
  .I0(sp_inst_32_dout[20]),
  .I1(sp_inst_33_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_621 (
  .O(mux_o_621),
  .I0(sp_inst_34_dout[20]),
  .I1(sp_inst_35_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_622 (
  .O(mux_o_622),
  .I0(sp_inst_36_dout[20]),
  .I1(sp_inst_37_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_623 (
  .O(mux_o_623),
  .I0(sp_inst_38_dout[20]),
  .I1(sp_inst_39_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_624 (
  .O(mux_o_624),
  .I0(sp_inst_40_dout[20]),
  .I1(sp_inst_41_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_625 (
  .O(mux_o_625),
  .I0(sp_inst_42_dout[20]),
  .I1(sp_inst_43_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_626 (
  .O(mux_o_626),
  .I0(sp_inst_44_dout[20]),
  .I1(sp_inst_45_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_627 (
  .O(mux_o_627),
  .I0(sp_inst_46_dout[20]),
  .I1(sp_inst_47_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_628 (
  .O(mux_o_628),
  .I0(sp_inst_48_dout[20]),
  .I1(sp_inst_49_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_629 (
  .O(mux_o_629),
  .I0(sp_inst_50_dout[20]),
  .I1(sp_inst_51_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_630 (
  .O(mux_o_630),
  .I0(sp_inst_52_dout[20]),
  .I1(sp_inst_53_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_631 (
  .O(mux_o_631),
  .I0(sp_inst_54_dout[20]),
  .I1(sp_inst_55_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_632 (
  .O(mux_o_632),
  .I0(sp_inst_56_dout[20]),
  .I1(sp_inst_57_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_633 (
  .O(mux_o_633),
  .I0(sp_inst_58_dout[20]),
  .I1(sp_inst_59_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_634 (
  .O(mux_o_634),
  .I0(sp_inst_60_dout[20]),
  .I1(sp_inst_61_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_635 (
  .O(mux_o_635),
  .I0(sp_inst_62_dout[20]),
  .I1(sp_inst_63_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_636 (
  .O(mux_o_636),
  .I0(mux_o_620),
  .I1(mux_o_621),
  .S0(dff_q_3)
);
MUX2 mux_inst_637 (
  .O(mux_o_637),
  .I0(mux_o_622),
  .I1(mux_o_623),
  .S0(dff_q_3)
);
MUX2 mux_inst_638 (
  .O(mux_o_638),
  .I0(mux_o_624),
  .I1(mux_o_625),
  .S0(dff_q_3)
);
MUX2 mux_inst_639 (
  .O(mux_o_639),
  .I0(mux_o_626),
  .I1(mux_o_627),
  .S0(dff_q_3)
);
MUX2 mux_inst_640 (
  .O(mux_o_640),
  .I0(mux_o_628),
  .I1(mux_o_629),
  .S0(dff_q_3)
);
MUX2 mux_inst_641 (
  .O(mux_o_641),
  .I0(mux_o_630),
  .I1(mux_o_631),
  .S0(dff_q_3)
);
MUX2 mux_inst_642 (
  .O(mux_o_642),
  .I0(mux_o_632),
  .I1(mux_o_633),
  .S0(dff_q_3)
);
MUX2 mux_inst_643 (
  .O(mux_o_643),
  .I0(mux_o_634),
  .I1(mux_o_635),
  .S0(dff_q_3)
);
MUX2 mux_inst_644 (
  .O(mux_o_644),
  .I0(mux_o_636),
  .I1(mux_o_637),
  .S0(dff_q_2)
);
MUX2 mux_inst_645 (
  .O(mux_o_645),
  .I0(mux_o_638),
  .I1(mux_o_639),
  .S0(dff_q_2)
);
MUX2 mux_inst_646 (
  .O(mux_o_646),
  .I0(mux_o_640),
  .I1(mux_o_641),
  .S0(dff_q_2)
);
MUX2 mux_inst_647 (
  .O(mux_o_647),
  .I0(mux_o_642),
  .I1(mux_o_643),
  .S0(dff_q_2)
);
MUX2 mux_inst_648 (
  .O(mux_o_648),
  .I0(mux_o_644),
  .I1(mux_o_645),
  .S0(dff_q_1)
);
MUX2 mux_inst_649 (
  .O(mux_o_649),
  .I0(mux_o_646),
  .I1(mux_o_647),
  .S0(dff_q_1)
);
MUX2 mux_inst_650 (
  .O(dout[20]),
  .I0(mux_o_648),
  .I1(mux_o_649),
  .S0(dff_q_0)
);
MUX2 mux_inst_651 (
  .O(mux_o_651),
  .I0(sp_inst_32_dout[21]),
  .I1(sp_inst_33_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_652 (
  .O(mux_o_652),
  .I0(sp_inst_34_dout[21]),
  .I1(sp_inst_35_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_653 (
  .O(mux_o_653),
  .I0(sp_inst_36_dout[21]),
  .I1(sp_inst_37_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_654 (
  .O(mux_o_654),
  .I0(sp_inst_38_dout[21]),
  .I1(sp_inst_39_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_655 (
  .O(mux_o_655),
  .I0(sp_inst_40_dout[21]),
  .I1(sp_inst_41_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_656 (
  .O(mux_o_656),
  .I0(sp_inst_42_dout[21]),
  .I1(sp_inst_43_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_657 (
  .O(mux_o_657),
  .I0(sp_inst_44_dout[21]),
  .I1(sp_inst_45_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_658 (
  .O(mux_o_658),
  .I0(sp_inst_46_dout[21]),
  .I1(sp_inst_47_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_659 (
  .O(mux_o_659),
  .I0(sp_inst_48_dout[21]),
  .I1(sp_inst_49_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_660 (
  .O(mux_o_660),
  .I0(sp_inst_50_dout[21]),
  .I1(sp_inst_51_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_661 (
  .O(mux_o_661),
  .I0(sp_inst_52_dout[21]),
  .I1(sp_inst_53_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_662 (
  .O(mux_o_662),
  .I0(sp_inst_54_dout[21]),
  .I1(sp_inst_55_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_663 (
  .O(mux_o_663),
  .I0(sp_inst_56_dout[21]),
  .I1(sp_inst_57_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_664 (
  .O(mux_o_664),
  .I0(sp_inst_58_dout[21]),
  .I1(sp_inst_59_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_665 (
  .O(mux_o_665),
  .I0(sp_inst_60_dout[21]),
  .I1(sp_inst_61_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_666 (
  .O(mux_o_666),
  .I0(sp_inst_62_dout[21]),
  .I1(sp_inst_63_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_667 (
  .O(mux_o_667),
  .I0(mux_o_651),
  .I1(mux_o_652),
  .S0(dff_q_3)
);
MUX2 mux_inst_668 (
  .O(mux_o_668),
  .I0(mux_o_653),
  .I1(mux_o_654),
  .S0(dff_q_3)
);
MUX2 mux_inst_669 (
  .O(mux_o_669),
  .I0(mux_o_655),
  .I1(mux_o_656),
  .S0(dff_q_3)
);
MUX2 mux_inst_670 (
  .O(mux_o_670),
  .I0(mux_o_657),
  .I1(mux_o_658),
  .S0(dff_q_3)
);
MUX2 mux_inst_671 (
  .O(mux_o_671),
  .I0(mux_o_659),
  .I1(mux_o_660),
  .S0(dff_q_3)
);
MUX2 mux_inst_672 (
  .O(mux_o_672),
  .I0(mux_o_661),
  .I1(mux_o_662),
  .S0(dff_q_3)
);
MUX2 mux_inst_673 (
  .O(mux_o_673),
  .I0(mux_o_663),
  .I1(mux_o_664),
  .S0(dff_q_3)
);
MUX2 mux_inst_674 (
  .O(mux_o_674),
  .I0(mux_o_665),
  .I1(mux_o_666),
  .S0(dff_q_3)
);
MUX2 mux_inst_675 (
  .O(mux_o_675),
  .I0(mux_o_667),
  .I1(mux_o_668),
  .S0(dff_q_2)
);
MUX2 mux_inst_676 (
  .O(mux_o_676),
  .I0(mux_o_669),
  .I1(mux_o_670),
  .S0(dff_q_2)
);
MUX2 mux_inst_677 (
  .O(mux_o_677),
  .I0(mux_o_671),
  .I1(mux_o_672),
  .S0(dff_q_2)
);
MUX2 mux_inst_678 (
  .O(mux_o_678),
  .I0(mux_o_673),
  .I1(mux_o_674),
  .S0(dff_q_2)
);
MUX2 mux_inst_679 (
  .O(mux_o_679),
  .I0(mux_o_675),
  .I1(mux_o_676),
  .S0(dff_q_1)
);
MUX2 mux_inst_680 (
  .O(mux_o_680),
  .I0(mux_o_677),
  .I1(mux_o_678),
  .S0(dff_q_1)
);
MUX2 mux_inst_681 (
  .O(dout[21]),
  .I0(mux_o_679),
  .I1(mux_o_680),
  .S0(dff_q_0)
);
MUX2 mux_inst_682 (
  .O(mux_o_682),
  .I0(sp_inst_32_dout[22]),
  .I1(sp_inst_33_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_683 (
  .O(mux_o_683),
  .I0(sp_inst_34_dout[22]),
  .I1(sp_inst_35_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_684 (
  .O(mux_o_684),
  .I0(sp_inst_36_dout[22]),
  .I1(sp_inst_37_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_685 (
  .O(mux_o_685),
  .I0(sp_inst_38_dout[22]),
  .I1(sp_inst_39_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_686 (
  .O(mux_o_686),
  .I0(sp_inst_40_dout[22]),
  .I1(sp_inst_41_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_687 (
  .O(mux_o_687),
  .I0(sp_inst_42_dout[22]),
  .I1(sp_inst_43_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_688 (
  .O(mux_o_688),
  .I0(sp_inst_44_dout[22]),
  .I1(sp_inst_45_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_689 (
  .O(mux_o_689),
  .I0(sp_inst_46_dout[22]),
  .I1(sp_inst_47_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_690 (
  .O(mux_o_690),
  .I0(sp_inst_48_dout[22]),
  .I1(sp_inst_49_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_691 (
  .O(mux_o_691),
  .I0(sp_inst_50_dout[22]),
  .I1(sp_inst_51_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_692 (
  .O(mux_o_692),
  .I0(sp_inst_52_dout[22]),
  .I1(sp_inst_53_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_693 (
  .O(mux_o_693),
  .I0(sp_inst_54_dout[22]),
  .I1(sp_inst_55_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_694 (
  .O(mux_o_694),
  .I0(sp_inst_56_dout[22]),
  .I1(sp_inst_57_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_695 (
  .O(mux_o_695),
  .I0(sp_inst_58_dout[22]),
  .I1(sp_inst_59_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_696 (
  .O(mux_o_696),
  .I0(sp_inst_60_dout[22]),
  .I1(sp_inst_61_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_697 (
  .O(mux_o_697),
  .I0(sp_inst_62_dout[22]),
  .I1(sp_inst_63_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_698 (
  .O(mux_o_698),
  .I0(mux_o_682),
  .I1(mux_o_683),
  .S0(dff_q_3)
);
MUX2 mux_inst_699 (
  .O(mux_o_699),
  .I0(mux_o_684),
  .I1(mux_o_685),
  .S0(dff_q_3)
);
MUX2 mux_inst_700 (
  .O(mux_o_700),
  .I0(mux_o_686),
  .I1(mux_o_687),
  .S0(dff_q_3)
);
MUX2 mux_inst_701 (
  .O(mux_o_701),
  .I0(mux_o_688),
  .I1(mux_o_689),
  .S0(dff_q_3)
);
MUX2 mux_inst_702 (
  .O(mux_o_702),
  .I0(mux_o_690),
  .I1(mux_o_691),
  .S0(dff_q_3)
);
MUX2 mux_inst_703 (
  .O(mux_o_703),
  .I0(mux_o_692),
  .I1(mux_o_693),
  .S0(dff_q_3)
);
MUX2 mux_inst_704 (
  .O(mux_o_704),
  .I0(mux_o_694),
  .I1(mux_o_695),
  .S0(dff_q_3)
);
MUX2 mux_inst_705 (
  .O(mux_o_705),
  .I0(mux_o_696),
  .I1(mux_o_697),
  .S0(dff_q_3)
);
MUX2 mux_inst_706 (
  .O(mux_o_706),
  .I0(mux_o_698),
  .I1(mux_o_699),
  .S0(dff_q_2)
);
MUX2 mux_inst_707 (
  .O(mux_o_707),
  .I0(mux_o_700),
  .I1(mux_o_701),
  .S0(dff_q_2)
);
MUX2 mux_inst_708 (
  .O(mux_o_708),
  .I0(mux_o_702),
  .I1(mux_o_703),
  .S0(dff_q_2)
);
MUX2 mux_inst_709 (
  .O(mux_o_709),
  .I0(mux_o_704),
  .I1(mux_o_705),
  .S0(dff_q_2)
);
MUX2 mux_inst_710 (
  .O(mux_o_710),
  .I0(mux_o_706),
  .I1(mux_o_707),
  .S0(dff_q_1)
);
MUX2 mux_inst_711 (
  .O(mux_o_711),
  .I0(mux_o_708),
  .I1(mux_o_709),
  .S0(dff_q_1)
);
MUX2 mux_inst_712 (
  .O(dout[22]),
  .I0(mux_o_710),
  .I1(mux_o_711),
  .S0(dff_q_0)
);
MUX2 mux_inst_713 (
  .O(mux_o_713),
  .I0(sp_inst_32_dout[23]),
  .I1(sp_inst_33_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_714 (
  .O(mux_o_714),
  .I0(sp_inst_34_dout[23]),
  .I1(sp_inst_35_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_715 (
  .O(mux_o_715),
  .I0(sp_inst_36_dout[23]),
  .I1(sp_inst_37_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_716 (
  .O(mux_o_716),
  .I0(sp_inst_38_dout[23]),
  .I1(sp_inst_39_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_717 (
  .O(mux_o_717),
  .I0(sp_inst_40_dout[23]),
  .I1(sp_inst_41_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_718 (
  .O(mux_o_718),
  .I0(sp_inst_42_dout[23]),
  .I1(sp_inst_43_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_719 (
  .O(mux_o_719),
  .I0(sp_inst_44_dout[23]),
  .I1(sp_inst_45_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_720 (
  .O(mux_o_720),
  .I0(sp_inst_46_dout[23]),
  .I1(sp_inst_47_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_721 (
  .O(mux_o_721),
  .I0(sp_inst_48_dout[23]),
  .I1(sp_inst_49_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_722 (
  .O(mux_o_722),
  .I0(sp_inst_50_dout[23]),
  .I1(sp_inst_51_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_723 (
  .O(mux_o_723),
  .I0(sp_inst_52_dout[23]),
  .I1(sp_inst_53_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_724 (
  .O(mux_o_724),
  .I0(sp_inst_54_dout[23]),
  .I1(sp_inst_55_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_725 (
  .O(mux_o_725),
  .I0(sp_inst_56_dout[23]),
  .I1(sp_inst_57_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_726 (
  .O(mux_o_726),
  .I0(sp_inst_58_dout[23]),
  .I1(sp_inst_59_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_727 (
  .O(mux_o_727),
  .I0(sp_inst_60_dout[23]),
  .I1(sp_inst_61_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_728 (
  .O(mux_o_728),
  .I0(sp_inst_62_dout[23]),
  .I1(sp_inst_63_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_729 (
  .O(mux_o_729),
  .I0(mux_o_713),
  .I1(mux_o_714),
  .S0(dff_q_3)
);
MUX2 mux_inst_730 (
  .O(mux_o_730),
  .I0(mux_o_715),
  .I1(mux_o_716),
  .S0(dff_q_3)
);
MUX2 mux_inst_731 (
  .O(mux_o_731),
  .I0(mux_o_717),
  .I1(mux_o_718),
  .S0(dff_q_3)
);
MUX2 mux_inst_732 (
  .O(mux_o_732),
  .I0(mux_o_719),
  .I1(mux_o_720),
  .S0(dff_q_3)
);
MUX2 mux_inst_733 (
  .O(mux_o_733),
  .I0(mux_o_721),
  .I1(mux_o_722),
  .S0(dff_q_3)
);
MUX2 mux_inst_734 (
  .O(mux_o_734),
  .I0(mux_o_723),
  .I1(mux_o_724),
  .S0(dff_q_3)
);
MUX2 mux_inst_735 (
  .O(mux_o_735),
  .I0(mux_o_725),
  .I1(mux_o_726),
  .S0(dff_q_3)
);
MUX2 mux_inst_736 (
  .O(mux_o_736),
  .I0(mux_o_727),
  .I1(mux_o_728),
  .S0(dff_q_3)
);
MUX2 mux_inst_737 (
  .O(mux_o_737),
  .I0(mux_o_729),
  .I1(mux_o_730),
  .S0(dff_q_2)
);
MUX2 mux_inst_738 (
  .O(mux_o_738),
  .I0(mux_o_731),
  .I1(mux_o_732),
  .S0(dff_q_2)
);
MUX2 mux_inst_739 (
  .O(mux_o_739),
  .I0(mux_o_733),
  .I1(mux_o_734),
  .S0(dff_q_2)
);
MUX2 mux_inst_740 (
  .O(mux_o_740),
  .I0(mux_o_735),
  .I1(mux_o_736),
  .S0(dff_q_2)
);
MUX2 mux_inst_741 (
  .O(mux_o_741),
  .I0(mux_o_737),
  .I1(mux_o_738),
  .S0(dff_q_1)
);
MUX2 mux_inst_742 (
  .O(mux_o_742),
  .I0(mux_o_739),
  .I1(mux_o_740),
  .S0(dff_q_1)
);
MUX2 mux_inst_743 (
  .O(dout[23]),
  .I0(mux_o_741),
  .I1(mux_o_742),
  .S0(dff_q_0)
);
MUX2 mux_inst_744 (
  .O(mux_o_744),
  .I0(sp_inst_32_dout[24]),
  .I1(sp_inst_33_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_745 (
  .O(mux_o_745),
  .I0(sp_inst_34_dout[24]),
  .I1(sp_inst_35_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_746 (
  .O(mux_o_746),
  .I0(sp_inst_36_dout[24]),
  .I1(sp_inst_37_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_747 (
  .O(mux_o_747),
  .I0(sp_inst_38_dout[24]),
  .I1(sp_inst_39_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_748 (
  .O(mux_o_748),
  .I0(sp_inst_40_dout[24]),
  .I1(sp_inst_41_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_749 (
  .O(mux_o_749),
  .I0(sp_inst_42_dout[24]),
  .I1(sp_inst_43_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_750 (
  .O(mux_o_750),
  .I0(sp_inst_44_dout[24]),
  .I1(sp_inst_45_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_751 (
  .O(mux_o_751),
  .I0(sp_inst_46_dout[24]),
  .I1(sp_inst_47_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_752 (
  .O(mux_o_752),
  .I0(sp_inst_48_dout[24]),
  .I1(sp_inst_49_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_753 (
  .O(mux_o_753),
  .I0(sp_inst_50_dout[24]),
  .I1(sp_inst_51_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_754 (
  .O(mux_o_754),
  .I0(sp_inst_52_dout[24]),
  .I1(sp_inst_53_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_755 (
  .O(mux_o_755),
  .I0(sp_inst_54_dout[24]),
  .I1(sp_inst_55_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_756 (
  .O(mux_o_756),
  .I0(sp_inst_56_dout[24]),
  .I1(sp_inst_57_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_757 (
  .O(mux_o_757),
  .I0(sp_inst_58_dout[24]),
  .I1(sp_inst_59_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_758 (
  .O(mux_o_758),
  .I0(sp_inst_60_dout[24]),
  .I1(sp_inst_61_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_759 (
  .O(mux_o_759),
  .I0(sp_inst_62_dout[24]),
  .I1(sp_inst_63_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_760 (
  .O(mux_o_760),
  .I0(mux_o_744),
  .I1(mux_o_745),
  .S0(dff_q_3)
);
MUX2 mux_inst_761 (
  .O(mux_o_761),
  .I0(mux_o_746),
  .I1(mux_o_747),
  .S0(dff_q_3)
);
MUX2 mux_inst_762 (
  .O(mux_o_762),
  .I0(mux_o_748),
  .I1(mux_o_749),
  .S0(dff_q_3)
);
MUX2 mux_inst_763 (
  .O(mux_o_763),
  .I0(mux_o_750),
  .I1(mux_o_751),
  .S0(dff_q_3)
);
MUX2 mux_inst_764 (
  .O(mux_o_764),
  .I0(mux_o_752),
  .I1(mux_o_753),
  .S0(dff_q_3)
);
MUX2 mux_inst_765 (
  .O(mux_o_765),
  .I0(mux_o_754),
  .I1(mux_o_755),
  .S0(dff_q_3)
);
MUX2 mux_inst_766 (
  .O(mux_o_766),
  .I0(mux_o_756),
  .I1(mux_o_757),
  .S0(dff_q_3)
);
MUX2 mux_inst_767 (
  .O(mux_o_767),
  .I0(mux_o_758),
  .I1(mux_o_759),
  .S0(dff_q_3)
);
MUX2 mux_inst_768 (
  .O(mux_o_768),
  .I0(mux_o_760),
  .I1(mux_o_761),
  .S0(dff_q_2)
);
MUX2 mux_inst_769 (
  .O(mux_o_769),
  .I0(mux_o_762),
  .I1(mux_o_763),
  .S0(dff_q_2)
);
MUX2 mux_inst_770 (
  .O(mux_o_770),
  .I0(mux_o_764),
  .I1(mux_o_765),
  .S0(dff_q_2)
);
MUX2 mux_inst_771 (
  .O(mux_o_771),
  .I0(mux_o_766),
  .I1(mux_o_767),
  .S0(dff_q_2)
);
MUX2 mux_inst_772 (
  .O(mux_o_772),
  .I0(mux_o_768),
  .I1(mux_o_769),
  .S0(dff_q_1)
);
MUX2 mux_inst_773 (
  .O(mux_o_773),
  .I0(mux_o_770),
  .I1(mux_o_771),
  .S0(dff_q_1)
);
MUX2 mux_inst_774 (
  .O(dout[24]),
  .I0(mux_o_772),
  .I1(mux_o_773),
  .S0(dff_q_0)
);
MUX2 mux_inst_775 (
  .O(mux_o_775),
  .I0(sp_inst_32_dout[25]),
  .I1(sp_inst_33_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_776 (
  .O(mux_o_776),
  .I0(sp_inst_34_dout[25]),
  .I1(sp_inst_35_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_777 (
  .O(mux_o_777),
  .I0(sp_inst_36_dout[25]),
  .I1(sp_inst_37_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_778 (
  .O(mux_o_778),
  .I0(sp_inst_38_dout[25]),
  .I1(sp_inst_39_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_779 (
  .O(mux_o_779),
  .I0(sp_inst_40_dout[25]),
  .I1(sp_inst_41_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_780 (
  .O(mux_o_780),
  .I0(sp_inst_42_dout[25]),
  .I1(sp_inst_43_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_781 (
  .O(mux_o_781),
  .I0(sp_inst_44_dout[25]),
  .I1(sp_inst_45_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_782 (
  .O(mux_o_782),
  .I0(sp_inst_46_dout[25]),
  .I1(sp_inst_47_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_783 (
  .O(mux_o_783),
  .I0(sp_inst_48_dout[25]),
  .I1(sp_inst_49_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_784 (
  .O(mux_o_784),
  .I0(sp_inst_50_dout[25]),
  .I1(sp_inst_51_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_785 (
  .O(mux_o_785),
  .I0(sp_inst_52_dout[25]),
  .I1(sp_inst_53_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_786 (
  .O(mux_o_786),
  .I0(sp_inst_54_dout[25]),
  .I1(sp_inst_55_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_787 (
  .O(mux_o_787),
  .I0(sp_inst_56_dout[25]),
  .I1(sp_inst_57_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_788 (
  .O(mux_o_788),
  .I0(sp_inst_58_dout[25]),
  .I1(sp_inst_59_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_789 (
  .O(mux_o_789),
  .I0(sp_inst_60_dout[25]),
  .I1(sp_inst_61_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_790 (
  .O(mux_o_790),
  .I0(sp_inst_62_dout[25]),
  .I1(sp_inst_63_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_791 (
  .O(mux_o_791),
  .I0(mux_o_775),
  .I1(mux_o_776),
  .S0(dff_q_3)
);
MUX2 mux_inst_792 (
  .O(mux_o_792),
  .I0(mux_o_777),
  .I1(mux_o_778),
  .S0(dff_q_3)
);
MUX2 mux_inst_793 (
  .O(mux_o_793),
  .I0(mux_o_779),
  .I1(mux_o_780),
  .S0(dff_q_3)
);
MUX2 mux_inst_794 (
  .O(mux_o_794),
  .I0(mux_o_781),
  .I1(mux_o_782),
  .S0(dff_q_3)
);
MUX2 mux_inst_795 (
  .O(mux_o_795),
  .I0(mux_o_783),
  .I1(mux_o_784),
  .S0(dff_q_3)
);
MUX2 mux_inst_796 (
  .O(mux_o_796),
  .I0(mux_o_785),
  .I1(mux_o_786),
  .S0(dff_q_3)
);
MUX2 mux_inst_797 (
  .O(mux_o_797),
  .I0(mux_o_787),
  .I1(mux_o_788),
  .S0(dff_q_3)
);
MUX2 mux_inst_798 (
  .O(mux_o_798),
  .I0(mux_o_789),
  .I1(mux_o_790),
  .S0(dff_q_3)
);
MUX2 mux_inst_799 (
  .O(mux_o_799),
  .I0(mux_o_791),
  .I1(mux_o_792),
  .S0(dff_q_2)
);
MUX2 mux_inst_800 (
  .O(mux_o_800),
  .I0(mux_o_793),
  .I1(mux_o_794),
  .S0(dff_q_2)
);
MUX2 mux_inst_801 (
  .O(mux_o_801),
  .I0(mux_o_795),
  .I1(mux_o_796),
  .S0(dff_q_2)
);
MUX2 mux_inst_802 (
  .O(mux_o_802),
  .I0(mux_o_797),
  .I1(mux_o_798),
  .S0(dff_q_2)
);
MUX2 mux_inst_803 (
  .O(mux_o_803),
  .I0(mux_o_799),
  .I1(mux_o_800),
  .S0(dff_q_1)
);
MUX2 mux_inst_804 (
  .O(mux_o_804),
  .I0(mux_o_801),
  .I1(mux_o_802),
  .S0(dff_q_1)
);
MUX2 mux_inst_805 (
  .O(dout[25]),
  .I0(mux_o_803),
  .I1(mux_o_804),
  .S0(dff_q_0)
);
MUX2 mux_inst_806 (
  .O(mux_o_806),
  .I0(sp_inst_32_dout[26]),
  .I1(sp_inst_33_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_807 (
  .O(mux_o_807),
  .I0(sp_inst_34_dout[26]),
  .I1(sp_inst_35_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_808 (
  .O(mux_o_808),
  .I0(sp_inst_36_dout[26]),
  .I1(sp_inst_37_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_809 (
  .O(mux_o_809),
  .I0(sp_inst_38_dout[26]),
  .I1(sp_inst_39_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_810 (
  .O(mux_o_810),
  .I0(sp_inst_40_dout[26]),
  .I1(sp_inst_41_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_811 (
  .O(mux_o_811),
  .I0(sp_inst_42_dout[26]),
  .I1(sp_inst_43_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_812 (
  .O(mux_o_812),
  .I0(sp_inst_44_dout[26]),
  .I1(sp_inst_45_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_813 (
  .O(mux_o_813),
  .I0(sp_inst_46_dout[26]),
  .I1(sp_inst_47_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_814 (
  .O(mux_o_814),
  .I0(sp_inst_48_dout[26]),
  .I1(sp_inst_49_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_815 (
  .O(mux_o_815),
  .I0(sp_inst_50_dout[26]),
  .I1(sp_inst_51_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_816 (
  .O(mux_o_816),
  .I0(sp_inst_52_dout[26]),
  .I1(sp_inst_53_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_817 (
  .O(mux_o_817),
  .I0(sp_inst_54_dout[26]),
  .I1(sp_inst_55_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_818 (
  .O(mux_o_818),
  .I0(sp_inst_56_dout[26]),
  .I1(sp_inst_57_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_819 (
  .O(mux_o_819),
  .I0(sp_inst_58_dout[26]),
  .I1(sp_inst_59_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_820 (
  .O(mux_o_820),
  .I0(sp_inst_60_dout[26]),
  .I1(sp_inst_61_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_821 (
  .O(mux_o_821),
  .I0(sp_inst_62_dout[26]),
  .I1(sp_inst_63_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_822 (
  .O(mux_o_822),
  .I0(mux_o_806),
  .I1(mux_o_807),
  .S0(dff_q_3)
);
MUX2 mux_inst_823 (
  .O(mux_o_823),
  .I0(mux_o_808),
  .I1(mux_o_809),
  .S0(dff_q_3)
);
MUX2 mux_inst_824 (
  .O(mux_o_824),
  .I0(mux_o_810),
  .I1(mux_o_811),
  .S0(dff_q_3)
);
MUX2 mux_inst_825 (
  .O(mux_o_825),
  .I0(mux_o_812),
  .I1(mux_o_813),
  .S0(dff_q_3)
);
MUX2 mux_inst_826 (
  .O(mux_o_826),
  .I0(mux_o_814),
  .I1(mux_o_815),
  .S0(dff_q_3)
);
MUX2 mux_inst_827 (
  .O(mux_o_827),
  .I0(mux_o_816),
  .I1(mux_o_817),
  .S0(dff_q_3)
);
MUX2 mux_inst_828 (
  .O(mux_o_828),
  .I0(mux_o_818),
  .I1(mux_o_819),
  .S0(dff_q_3)
);
MUX2 mux_inst_829 (
  .O(mux_o_829),
  .I0(mux_o_820),
  .I1(mux_o_821),
  .S0(dff_q_3)
);
MUX2 mux_inst_830 (
  .O(mux_o_830),
  .I0(mux_o_822),
  .I1(mux_o_823),
  .S0(dff_q_2)
);
MUX2 mux_inst_831 (
  .O(mux_o_831),
  .I0(mux_o_824),
  .I1(mux_o_825),
  .S0(dff_q_2)
);
MUX2 mux_inst_832 (
  .O(mux_o_832),
  .I0(mux_o_826),
  .I1(mux_o_827),
  .S0(dff_q_2)
);
MUX2 mux_inst_833 (
  .O(mux_o_833),
  .I0(mux_o_828),
  .I1(mux_o_829),
  .S0(dff_q_2)
);
MUX2 mux_inst_834 (
  .O(mux_o_834),
  .I0(mux_o_830),
  .I1(mux_o_831),
  .S0(dff_q_1)
);
MUX2 mux_inst_835 (
  .O(mux_o_835),
  .I0(mux_o_832),
  .I1(mux_o_833),
  .S0(dff_q_1)
);
MUX2 mux_inst_836 (
  .O(dout[26]),
  .I0(mux_o_834),
  .I1(mux_o_835),
  .S0(dff_q_0)
);
MUX2 mux_inst_837 (
  .O(mux_o_837),
  .I0(sp_inst_32_dout[27]),
  .I1(sp_inst_33_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_838 (
  .O(mux_o_838),
  .I0(sp_inst_34_dout[27]),
  .I1(sp_inst_35_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_839 (
  .O(mux_o_839),
  .I0(sp_inst_36_dout[27]),
  .I1(sp_inst_37_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_840 (
  .O(mux_o_840),
  .I0(sp_inst_38_dout[27]),
  .I1(sp_inst_39_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_841 (
  .O(mux_o_841),
  .I0(sp_inst_40_dout[27]),
  .I1(sp_inst_41_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_842 (
  .O(mux_o_842),
  .I0(sp_inst_42_dout[27]),
  .I1(sp_inst_43_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_843 (
  .O(mux_o_843),
  .I0(sp_inst_44_dout[27]),
  .I1(sp_inst_45_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_844 (
  .O(mux_o_844),
  .I0(sp_inst_46_dout[27]),
  .I1(sp_inst_47_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_845 (
  .O(mux_o_845),
  .I0(sp_inst_48_dout[27]),
  .I1(sp_inst_49_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_846 (
  .O(mux_o_846),
  .I0(sp_inst_50_dout[27]),
  .I1(sp_inst_51_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_847 (
  .O(mux_o_847),
  .I0(sp_inst_52_dout[27]),
  .I1(sp_inst_53_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_848 (
  .O(mux_o_848),
  .I0(sp_inst_54_dout[27]),
  .I1(sp_inst_55_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_849 (
  .O(mux_o_849),
  .I0(sp_inst_56_dout[27]),
  .I1(sp_inst_57_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_850 (
  .O(mux_o_850),
  .I0(sp_inst_58_dout[27]),
  .I1(sp_inst_59_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_851 (
  .O(mux_o_851),
  .I0(sp_inst_60_dout[27]),
  .I1(sp_inst_61_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_852 (
  .O(mux_o_852),
  .I0(sp_inst_62_dout[27]),
  .I1(sp_inst_63_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_853 (
  .O(mux_o_853),
  .I0(mux_o_837),
  .I1(mux_o_838),
  .S0(dff_q_3)
);
MUX2 mux_inst_854 (
  .O(mux_o_854),
  .I0(mux_o_839),
  .I1(mux_o_840),
  .S0(dff_q_3)
);
MUX2 mux_inst_855 (
  .O(mux_o_855),
  .I0(mux_o_841),
  .I1(mux_o_842),
  .S0(dff_q_3)
);
MUX2 mux_inst_856 (
  .O(mux_o_856),
  .I0(mux_o_843),
  .I1(mux_o_844),
  .S0(dff_q_3)
);
MUX2 mux_inst_857 (
  .O(mux_o_857),
  .I0(mux_o_845),
  .I1(mux_o_846),
  .S0(dff_q_3)
);
MUX2 mux_inst_858 (
  .O(mux_o_858),
  .I0(mux_o_847),
  .I1(mux_o_848),
  .S0(dff_q_3)
);
MUX2 mux_inst_859 (
  .O(mux_o_859),
  .I0(mux_o_849),
  .I1(mux_o_850),
  .S0(dff_q_3)
);
MUX2 mux_inst_860 (
  .O(mux_o_860),
  .I0(mux_o_851),
  .I1(mux_o_852),
  .S0(dff_q_3)
);
MUX2 mux_inst_861 (
  .O(mux_o_861),
  .I0(mux_o_853),
  .I1(mux_o_854),
  .S0(dff_q_2)
);
MUX2 mux_inst_862 (
  .O(mux_o_862),
  .I0(mux_o_855),
  .I1(mux_o_856),
  .S0(dff_q_2)
);
MUX2 mux_inst_863 (
  .O(mux_o_863),
  .I0(mux_o_857),
  .I1(mux_o_858),
  .S0(dff_q_2)
);
MUX2 mux_inst_864 (
  .O(mux_o_864),
  .I0(mux_o_859),
  .I1(mux_o_860),
  .S0(dff_q_2)
);
MUX2 mux_inst_865 (
  .O(mux_o_865),
  .I0(mux_o_861),
  .I1(mux_o_862),
  .S0(dff_q_1)
);
MUX2 mux_inst_866 (
  .O(mux_o_866),
  .I0(mux_o_863),
  .I1(mux_o_864),
  .S0(dff_q_1)
);
MUX2 mux_inst_867 (
  .O(dout[27]),
  .I0(mux_o_865),
  .I1(mux_o_866),
  .S0(dff_q_0)
);
MUX2 mux_inst_868 (
  .O(mux_o_868),
  .I0(sp_inst_32_dout[28]),
  .I1(sp_inst_33_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_869 (
  .O(mux_o_869),
  .I0(sp_inst_34_dout[28]),
  .I1(sp_inst_35_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_870 (
  .O(mux_o_870),
  .I0(sp_inst_36_dout[28]),
  .I1(sp_inst_37_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_871 (
  .O(mux_o_871),
  .I0(sp_inst_38_dout[28]),
  .I1(sp_inst_39_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_872 (
  .O(mux_o_872),
  .I0(sp_inst_40_dout[28]),
  .I1(sp_inst_41_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_873 (
  .O(mux_o_873),
  .I0(sp_inst_42_dout[28]),
  .I1(sp_inst_43_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_874 (
  .O(mux_o_874),
  .I0(sp_inst_44_dout[28]),
  .I1(sp_inst_45_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_875 (
  .O(mux_o_875),
  .I0(sp_inst_46_dout[28]),
  .I1(sp_inst_47_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_876 (
  .O(mux_o_876),
  .I0(sp_inst_48_dout[28]),
  .I1(sp_inst_49_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_877 (
  .O(mux_o_877),
  .I0(sp_inst_50_dout[28]),
  .I1(sp_inst_51_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_878 (
  .O(mux_o_878),
  .I0(sp_inst_52_dout[28]),
  .I1(sp_inst_53_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_879 (
  .O(mux_o_879),
  .I0(sp_inst_54_dout[28]),
  .I1(sp_inst_55_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_880 (
  .O(mux_o_880),
  .I0(sp_inst_56_dout[28]),
  .I1(sp_inst_57_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_881 (
  .O(mux_o_881),
  .I0(sp_inst_58_dout[28]),
  .I1(sp_inst_59_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_882 (
  .O(mux_o_882),
  .I0(sp_inst_60_dout[28]),
  .I1(sp_inst_61_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_883 (
  .O(mux_o_883),
  .I0(sp_inst_62_dout[28]),
  .I1(sp_inst_63_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_884 (
  .O(mux_o_884),
  .I0(mux_o_868),
  .I1(mux_o_869),
  .S0(dff_q_3)
);
MUX2 mux_inst_885 (
  .O(mux_o_885),
  .I0(mux_o_870),
  .I1(mux_o_871),
  .S0(dff_q_3)
);
MUX2 mux_inst_886 (
  .O(mux_o_886),
  .I0(mux_o_872),
  .I1(mux_o_873),
  .S0(dff_q_3)
);
MUX2 mux_inst_887 (
  .O(mux_o_887),
  .I0(mux_o_874),
  .I1(mux_o_875),
  .S0(dff_q_3)
);
MUX2 mux_inst_888 (
  .O(mux_o_888),
  .I0(mux_o_876),
  .I1(mux_o_877),
  .S0(dff_q_3)
);
MUX2 mux_inst_889 (
  .O(mux_o_889),
  .I0(mux_o_878),
  .I1(mux_o_879),
  .S0(dff_q_3)
);
MUX2 mux_inst_890 (
  .O(mux_o_890),
  .I0(mux_o_880),
  .I1(mux_o_881),
  .S0(dff_q_3)
);
MUX2 mux_inst_891 (
  .O(mux_o_891),
  .I0(mux_o_882),
  .I1(mux_o_883),
  .S0(dff_q_3)
);
MUX2 mux_inst_892 (
  .O(mux_o_892),
  .I0(mux_o_884),
  .I1(mux_o_885),
  .S0(dff_q_2)
);
MUX2 mux_inst_893 (
  .O(mux_o_893),
  .I0(mux_o_886),
  .I1(mux_o_887),
  .S0(dff_q_2)
);
MUX2 mux_inst_894 (
  .O(mux_o_894),
  .I0(mux_o_888),
  .I1(mux_o_889),
  .S0(dff_q_2)
);
MUX2 mux_inst_895 (
  .O(mux_o_895),
  .I0(mux_o_890),
  .I1(mux_o_891),
  .S0(dff_q_2)
);
MUX2 mux_inst_896 (
  .O(mux_o_896),
  .I0(mux_o_892),
  .I1(mux_o_893),
  .S0(dff_q_1)
);
MUX2 mux_inst_897 (
  .O(mux_o_897),
  .I0(mux_o_894),
  .I1(mux_o_895),
  .S0(dff_q_1)
);
MUX2 mux_inst_898 (
  .O(dout[28]),
  .I0(mux_o_896),
  .I1(mux_o_897),
  .S0(dff_q_0)
);
MUX2 mux_inst_899 (
  .O(mux_o_899),
  .I0(sp_inst_32_dout[29]),
  .I1(sp_inst_33_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_900 (
  .O(mux_o_900),
  .I0(sp_inst_34_dout[29]),
  .I1(sp_inst_35_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_901 (
  .O(mux_o_901),
  .I0(sp_inst_36_dout[29]),
  .I1(sp_inst_37_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_902 (
  .O(mux_o_902),
  .I0(sp_inst_38_dout[29]),
  .I1(sp_inst_39_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_903 (
  .O(mux_o_903),
  .I0(sp_inst_40_dout[29]),
  .I1(sp_inst_41_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_904 (
  .O(mux_o_904),
  .I0(sp_inst_42_dout[29]),
  .I1(sp_inst_43_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_905 (
  .O(mux_o_905),
  .I0(sp_inst_44_dout[29]),
  .I1(sp_inst_45_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_906 (
  .O(mux_o_906),
  .I0(sp_inst_46_dout[29]),
  .I1(sp_inst_47_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_907 (
  .O(mux_o_907),
  .I0(sp_inst_48_dout[29]),
  .I1(sp_inst_49_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_908 (
  .O(mux_o_908),
  .I0(sp_inst_50_dout[29]),
  .I1(sp_inst_51_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_909 (
  .O(mux_o_909),
  .I0(sp_inst_52_dout[29]),
  .I1(sp_inst_53_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_910 (
  .O(mux_o_910),
  .I0(sp_inst_54_dout[29]),
  .I1(sp_inst_55_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_911 (
  .O(mux_o_911),
  .I0(sp_inst_56_dout[29]),
  .I1(sp_inst_57_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_912 (
  .O(mux_o_912),
  .I0(sp_inst_58_dout[29]),
  .I1(sp_inst_59_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_913 (
  .O(mux_o_913),
  .I0(sp_inst_60_dout[29]),
  .I1(sp_inst_61_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_914 (
  .O(mux_o_914),
  .I0(sp_inst_62_dout[29]),
  .I1(sp_inst_63_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_915 (
  .O(mux_o_915),
  .I0(mux_o_899),
  .I1(mux_o_900),
  .S0(dff_q_3)
);
MUX2 mux_inst_916 (
  .O(mux_o_916),
  .I0(mux_o_901),
  .I1(mux_o_902),
  .S0(dff_q_3)
);
MUX2 mux_inst_917 (
  .O(mux_o_917),
  .I0(mux_o_903),
  .I1(mux_o_904),
  .S0(dff_q_3)
);
MUX2 mux_inst_918 (
  .O(mux_o_918),
  .I0(mux_o_905),
  .I1(mux_o_906),
  .S0(dff_q_3)
);
MUX2 mux_inst_919 (
  .O(mux_o_919),
  .I0(mux_o_907),
  .I1(mux_o_908),
  .S0(dff_q_3)
);
MUX2 mux_inst_920 (
  .O(mux_o_920),
  .I0(mux_o_909),
  .I1(mux_o_910),
  .S0(dff_q_3)
);
MUX2 mux_inst_921 (
  .O(mux_o_921),
  .I0(mux_o_911),
  .I1(mux_o_912),
  .S0(dff_q_3)
);
MUX2 mux_inst_922 (
  .O(mux_o_922),
  .I0(mux_o_913),
  .I1(mux_o_914),
  .S0(dff_q_3)
);
MUX2 mux_inst_923 (
  .O(mux_o_923),
  .I0(mux_o_915),
  .I1(mux_o_916),
  .S0(dff_q_2)
);
MUX2 mux_inst_924 (
  .O(mux_o_924),
  .I0(mux_o_917),
  .I1(mux_o_918),
  .S0(dff_q_2)
);
MUX2 mux_inst_925 (
  .O(mux_o_925),
  .I0(mux_o_919),
  .I1(mux_o_920),
  .S0(dff_q_2)
);
MUX2 mux_inst_926 (
  .O(mux_o_926),
  .I0(mux_o_921),
  .I1(mux_o_922),
  .S0(dff_q_2)
);
MUX2 mux_inst_927 (
  .O(mux_o_927),
  .I0(mux_o_923),
  .I1(mux_o_924),
  .S0(dff_q_1)
);
MUX2 mux_inst_928 (
  .O(mux_o_928),
  .I0(mux_o_925),
  .I1(mux_o_926),
  .S0(dff_q_1)
);
MUX2 mux_inst_929 (
  .O(dout[29]),
  .I0(mux_o_927),
  .I1(mux_o_928),
  .S0(dff_q_0)
);
MUX2 mux_inst_930 (
  .O(mux_o_930),
  .I0(sp_inst_32_dout[30]),
  .I1(sp_inst_33_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_931 (
  .O(mux_o_931),
  .I0(sp_inst_34_dout[30]),
  .I1(sp_inst_35_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_932 (
  .O(mux_o_932),
  .I0(sp_inst_36_dout[30]),
  .I1(sp_inst_37_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_933 (
  .O(mux_o_933),
  .I0(sp_inst_38_dout[30]),
  .I1(sp_inst_39_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_934 (
  .O(mux_o_934),
  .I0(sp_inst_40_dout[30]),
  .I1(sp_inst_41_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_935 (
  .O(mux_o_935),
  .I0(sp_inst_42_dout[30]),
  .I1(sp_inst_43_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_936 (
  .O(mux_o_936),
  .I0(sp_inst_44_dout[30]),
  .I1(sp_inst_45_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_937 (
  .O(mux_o_937),
  .I0(sp_inst_46_dout[30]),
  .I1(sp_inst_47_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_938 (
  .O(mux_o_938),
  .I0(sp_inst_48_dout[30]),
  .I1(sp_inst_49_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_939 (
  .O(mux_o_939),
  .I0(sp_inst_50_dout[30]),
  .I1(sp_inst_51_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_940 (
  .O(mux_o_940),
  .I0(sp_inst_52_dout[30]),
  .I1(sp_inst_53_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_941 (
  .O(mux_o_941),
  .I0(sp_inst_54_dout[30]),
  .I1(sp_inst_55_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_942 (
  .O(mux_o_942),
  .I0(sp_inst_56_dout[30]),
  .I1(sp_inst_57_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_943 (
  .O(mux_o_943),
  .I0(sp_inst_58_dout[30]),
  .I1(sp_inst_59_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_944 (
  .O(mux_o_944),
  .I0(sp_inst_60_dout[30]),
  .I1(sp_inst_61_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_945 (
  .O(mux_o_945),
  .I0(sp_inst_62_dout[30]),
  .I1(sp_inst_63_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_946 (
  .O(mux_o_946),
  .I0(mux_o_930),
  .I1(mux_o_931),
  .S0(dff_q_3)
);
MUX2 mux_inst_947 (
  .O(mux_o_947),
  .I0(mux_o_932),
  .I1(mux_o_933),
  .S0(dff_q_3)
);
MUX2 mux_inst_948 (
  .O(mux_o_948),
  .I0(mux_o_934),
  .I1(mux_o_935),
  .S0(dff_q_3)
);
MUX2 mux_inst_949 (
  .O(mux_o_949),
  .I0(mux_o_936),
  .I1(mux_o_937),
  .S0(dff_q_3)
);
MUX2 mux_inst_950 (
  .O(mux_o_950),
  .I0(mux_o_938),
  .I1(mux_o_939),
  .S0(dff_q_3)
);
MUX2 mux_inst_951 (
  .O(mux_o_951),
  .I0(mux_o_940),
  .I1(mux_o_941),
  .S0(dff_q_3)
);
MUX2 mux_inst_952 (
  .O(mux_o_952),
  .I0(mux_o_942),
  .I1(mux_o_943),
  .S0(dff_q_3)
);
MUX2 mux_inst_953 (
  .O(mux_o_953),
  .I0(mux_o_944),
  .I1(mux_o_945),
  .S0(dff_q_3)
);
MUX2 mux_inst_954 (
  .O(mux_o_954),
  .I0(mux_o_946),
  .I1(mux_o_947),
  .S0(dff_q_2)
);
MUX2 mux_inst_955 (
  .O(mux_o_955),
  .I0(mux_o_948),
  .I1(mux_o_949),
  .S0(dff_q_2)
);
MUX2 mux_inst_956 (
  .O(mux_o_956),
  .I0(mux_o_950),
  .I1(mux_o_951),
  .S0(dff_q_2)
);
MUX2 mux_inst_957 (
  .O(mux_o_957),
  .I0(mux_o_952),
  .I1(mux_o_953),
  .S0(dff_q_2)
);
MUX2 mux_inst_958 (
  .O(mux_o_958),
  .I0(mux_o_954),
  .I1(mux_o_955),
  .S0(dff_q_1)
);
MUX2 mux_inst_959 (
  .O(mux_o_959),
  .I0(mux_o_956),
  .I1(mux_o_957),
  .S0(dff_q_1)
);
MUX2 mux_inst_960 (
  .O(dout[30]),
  .I0(mux_o_958),
  .I1(mux_o_959),
  .S0(dff_q_0)
);
MUX2 mux_inst_961 (
  .O(mux_o_961),
  .I0(sp_inst_32_dout[31]),
  .I1(sp_inst_33_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_962 (
  .O(mux_o_962),
  .I0(sp_inst_34_dout[31]),
  .I1(sp_inst_35_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_963 (
  .O(mux_o_963),
  .I0(sp_inst_36_dout[31]),
  .I1(sp_inst_37_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_964 (
  .O(mux_o_964),
  .I0(sp_inst_38_dout[31]),
  .I1(sp_inst_39_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_965 (
  .O(mux_o_965),
  .I0(sp_inst_40_dout[31]),
  .I1(sp_inst_41_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_966 (
  .O(mux_o_966),
  .I0(sp_inst_42_dout[31]),
  .I1(sp_inst_43_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_967 (
  .O(mux_o_967),
  .I0(sp_inst_44_dout[31]),
  .I1(sp_inst_45_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_968 (
  .O(mux_o_968),
  .I0(sp_inst_46_dout[31]),
  .I1(sp_inst_47_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_969 (
  .O(mux_o_969),
  .I0(sp_inst_48_dout[31]),
  .I1(sp_inst_49_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_970 (
  .O(mux_o_970),
  .I0(sp_inst_50_dout[31]),
  .I1(sp_inst_51_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_971 (
  .O(mux_o_971),
  .I0(sp_inst_52_dout[31]),
  .I1(sp_inst_53_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_972 (
  .O(mux_o_972),
  .I0(sp_inst_54_dout[31]),
  .I1(sp_inst_55_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_973 (
  .O(mux_o_973),
  .I0(sp_inst_56_dout[31]),
  .I1(sp_inst_57_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_974 (
  .O(mux_o_974),
  .I0(sp_inst_58_dout[31]),
  .I1(sp_inst_59_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_975 (
  .O(mux_o_975),
  .I0(sp_inst_60_dout[31]),
  .I1(sp_inst_61_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_976 (
  .O(mux_o_976),
  .I0(sp_inst_62_dout[31]),
  .I1(sp_inst_63_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_977 (
  .O(mux_o_977),
  .I0(mux_o_961),
  .I1(mux_o_962),
  .S0(dff_q_3)
);
MUX2 mux_inst_978 (
  .O(mux_o_978),
  .I0(mux_o_963),
  .I1(mux_o_964),
  .S0(dff_q_3)
);
MUX2 mux_inst_979 (
  .O(mux_o_979),
  .I0(mux_o_965),
  .I1(mux_o_966),
  .S0(dff_q_3)
);
MUX2 mux_inst_980 (
  .O(mux_o_980),
  .I0(mux_o_967),
  .I1(mux_o_968),
  .S0(dff_q_3)
);
MUX2 mux_inst_981 (
  .O(mux_o_981),
  .I0(mux_o_969),
  .I1(mux_o_970),
  .S0(dff_q_3)
);
MUX2 mux_inst_982 (
  .O(mux_o_982),
  .I0(mux_o_971),
  .I1(mux_o_972),
  .S0(dff_q_3)
);
MUX2 mux_inst_983 (
  .O(mux_o_983),
  .I0(mux_o_973),
  .I1(mux_o_974),
  .S0(dff_q_3)
);
MUX2 mux_inst_984 (
  .O(mux_o_984),
  .I0(mux_o_975),
  .I1(mux_o_976),
  .S0(dff_q_3)
);
MUX2 mux_inst_985 (
  .O(mux_o_985),
  .I0(mux_o_977),
  .I1(mux_o_978),
  .S0(dff_q_2)
);
MUX2 mux_inst_986 (
  .O(mux_o_986),
  .I0(mux_o_979),
  .I1(mux_o_980),
  .S0(dff_q_2)
);
MUX2 mux_inst_987 (
  .O(mux_o_987),
  .I0(mux_o_981),
  .I1(mux_o_982),
  .S0(dff_q_2)
);
MUX2 mux_inst_988 (
  .O(mux_o_988),
  .I0(mux_o_983),
  .I1(mux_o_984),
  .S0(dff_q_2)
);
MUX2 mux_inst_989 (
  .O(mux_o_989),
  .I0(mux_o_985),
  .I1(mux_o_986),
  .S0(dff_q_1)
);
MUX2 mux_inst_990 (
  .O(mux_o_990),
  .I0(mux_o_987),
  .I1(mux_o_988),
  .S0(dff_q_1)
);
MUX2 mux_inst_991 (
  .O(dout[31]),
  .I0(mux_o_989),
  .I1(mux_o_990),
  .S0(dff_q_0)
);
endmodule //Gowin_SP
