//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.01 (64-bit)
//Part Number: GW5AST-LV138FPG676AES
//Device: GW5AST-138B
//Device Version: B
//Created Time: Fri Apr 19 21:29:28 2024

module blk_mem_gen_0 (dout, clk, oce, ce, reset, wre, ad, din, byte_en);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [14:0] ad;
input [31:0] din;
input [3:0] byte_en;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire [15:0] sp_inst_0_dout_w;
wire [15:0] sp_inst_0_dout;
wire [15:0] sp_inst_1_dout_w;
wire [15:0] sp_inst_1_dout;
wire [15:0] sp_inst_2_dout_w;
wire [15:0] sp_inst_2_dout;
wire [15:0] sp_inst_3_dout_w;
wire [15:0] sp_inst_3_dout;
wire [15:0] sp_inst_4_dout_w;
wire [15:0] sp_inst_4_dout;
wire [15:0] sp_inst_5_dout_w;
wire [15:0] sp_inst_5_dout;
wire [15:0] sp_inst_6_dout_w;
wire [15:0] sp_inst_6_dout;
wire [15:0] sp_inst_7_dout_w;
wire [15:0] sp_inst_7_dout;
wire [15:0] sp_inst_8_dout_w;
wire [15:0] sp_inst_8_dout;
wire [15:0] sp_inst_9_dout_w;
wire [15:0] sp_inst_9_dout;
wire [15:0] sp_inst_10_dout_w;
wire [15:0] sp_inst_10_dout;
wire [15:0] sp_inst_11_dout_w;
wire [15:0] sp_inst_11_dout;
wire [15:0] sp_inst_12_dout_w;
wire [15:0] sp_inst_12_dout;
wire [15:0] sp_inst_13_dout_w;
wire [15:0] sp_inst_13_dout;
wire [15:0] sp_inst_14_dout_w;
wire [15:0] sp_inst_14_dout;
wire [15:0] sp_inst_15_dout_w;
wire [15:0] sp_inst_15_dout;
wire [15:0] sp_inst_16_dout_w;
wire [15:0] sp_inst_16_dout;
wire [15:0] sp_inst_17_dout_w;
wire [15:0] sp_inst_17_dout;
wire [15:0] sp_inst_18_dout_w;
wire [15:0] sp_inst_18_dout;
wire [15:0] sp_inst_19_dout_w;
wire [15:0] sp_inst_19_dout;
wire [15:0] sp_inst_20_dout_w;
wire [15:0] sp_inst_20_dout;
wire [15:0] sp_inst_21_dout_w;
wire [15:0] sp_inst_21_dout;
wire [15:0] sp_inst_22_dout_w;
wire [15:0] sp_inst_22_dout;
wire [15:0] sp_inst_23_dout_w;
wire [15:0] sp_inst_23_dout;
wire [15:0] sp_inst_24_dout_w;
wire [15:0] sp_inst_24_dout;
wire [15:0] sp_inst_25_dout_w;
wire [15:0] sp_inst_25_dout;
wire [15:0] sp_inst_26_dout_w;
wire [15:0] sp_inst_26_dout;
wire [15:0] sp_inst_27_dout_w;
wire [15:0] sp_inst_27_dout;
wire [15:0] sp_inst_28_dout_w;
wire [15:0] sp_inst_28_dout;
wire [15:0] sp_inst_29_dout_w;
wire [15:0] sp_inst_29_dout;
wire [15:0] sp_inst_30_dout_w;
wire [15:0] sp_inst_30_dout;
wire [15:0] sp_inst_31_dout_w;
wire [15:0] sp_inst_31_dout;
wire [15:0] sp_inst_32_dout_w;
wire [31:16] sp_inst_32_dout;
wire [15:0] sp_inst_33_dout_w;
wire [31:16] sp_inst_33_dout;
wire [15:0] sp_inst_34_dout_w;
wire [31:16] sp_inst_34_dout;
wire [15:0] sp_inst_35_dout_w;
wire [31:16] sp_inst_35_dout;
wire [15:0] sp_inst_36_dout_w;
wire [31:16] sp_inst_36_dout;
wire [15:0] sp_inst_37_dout_w;
wire [31:16] sp_inst_37_dout;
wire [15:0] sp_inst_38_dout_w;
wire [31:16] sp_inst_38_dout;
wire [15:0] sp_inst_39_dout_w;
wire [31:16] sp_inst_39_dout;
wire [15:0] sp_inst_40_dout_w;
wire [31:16] sp_inst_40_dout;
wire [15:0] sp_inst_41_dout_w;
wire [31:16] sp_inst_41_dout;
wire [15:0] sp_inst_42_dout_w;
wire [31:16] sp_inst_42_dout;
wire [15:0] sp_inst_43_dout_w;
wire [31:16] sp_inst_43_dout;
wire [15:0] sp_inst_44_dout_w;
wire [31:16] sp_inst_44_dout;
wire [15:0] sp_inst_45_dout_w;
wire [31:16] sp_inst_45_dout;
wire [15:0] sp_inst_46_dout_w;
wire [31:16] sp_inst_46_dout;
wire [15:0] sp_inst_47_dout_w;
wire [31:16] sp_inst_47_dout;
wire [15:0] sp_inst_48_dout_w;
wire [31:16] sp_inst_48_dout;
wire [15:0] sp_inst_49_dout_w;
wire [31:16] sp_inst_49_dout;
wire [15:0] sp_inst_50_dout_w;
wire [31:16] sp_inst_50_dout;
wire [15:0] sp_inst_51_dout_w;
wire [31:16] sp_inst_51_dout;
wire [15:0] sp_inst_52_dout_w;
wire [31:16] sp_inst_52_dout;
wire [15:0] sp_inst_53_dout_w;
wire [31:16] sp_inst_53_dout;
wire [15:0] sp_inst_54_dout_w;
wire [31:16] sp_inst_54_dout;
wire [15:0] sp_inst_55_dout_w;
wire [31:16] sp_inst_55_dout;
wire [15:0] sp_inst_56_dout_w;
wire [31:16] sp_inst_56_dout;
wire [15:0] sp_inst_57_dout_w;
wire [31:16] sp_inst_57_dout;
wire [15:0] sp_inst_58_dout_w;
wire [31:16] sp_inst_58_dout;
wire [15:0] sp_inst_59_dout_w;
wire [31:16] sp_inst_59_dout;
wire [15:0] sp_inst_60_dout_w;
wire [31:16] sp_inst_60_dout;
wire [15:0] sp_inst_61_dout_w;
wire [31:16] sp_inst_61_dout;
wire [15:0] sp_inst_62_dout_w;
wire [31:16] sp_inst_62_dout;
wire [15:0] sp_inst_63_dout_w;
wire [31:16] sp_inst_63_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_91;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_104;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_124;
wire mux_o_125;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_164;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_179;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_209;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_224;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_245;
wire mux_o_246;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_251;
wire mux_o_252;
wire mux_o_253;
wire mux_o_254;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_258;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_265;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_269;
wire mux_o_270;
wire mux_o_271;
wire mux_o_272;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_279;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_284;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_299;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_308;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_314;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_321;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_329;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_335;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_349;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_356;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_360;
wire mux_o_361;
wire mux_o_362;
wire mux_o_363;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_370;
wire mux_o_372;
wire mux_o_373;
wire mux_o_374;
wire mux_o_375;
wire mux_o_376;
wire mux_o_377;
wire mux_o_378;
wire mux_o_379;
wire mux_o_380;
wire mux_o_381;
wire mux_o_382;
wire mux_o_383;
wire mux_o_384;
wire mux_o_385;
wire mux_o_386;
wire mux_o_387;
wire mux_o_388;
wire mux_o_389;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_401;
wire mux_o_403;
wire mux_o_404;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_408;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_412;
wire mux_o_413;
wire mux_o_414;
wire mux_o_415;
wire mux_o_416;
wire mux_o_417;
wire mux_o_418;
wire mux_o_419;
wire mux_o_420;
wire mux_o_421;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_426;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_431;
wire mux_o_432;
wire mux_o_434;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_440;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_449;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_453;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_460;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_465;
wire mux_o_466;
wire mux_o_467;
wire mux_o_468;
wire mux_o_469;
wire mux_o_470;
wire mux_o_471;
wire mux_o_472;
wire mux_o_473;
wire mux_o_474;
wire mux_o_475;
wire mux_o_476;
wire mux_o_477;
wire mux_o_478;
wire mux_o_479;
wire mux_o_480;
wire mux_o_481;
wire mux_o_482;
wire mux_o_483;
wire mux_o_484;
wire mux_o_485;
wire mux_o_486;
wire mux_o_487;
wire mux_o_488;
wire mux_o_489;
wire mux_o_490;
wire mux_o_491;
wire mux_o_492;
wire mux_o_493;
wire mux_o_494;
wire mux_o_496;
wire mux_o_497;
wire mux_o_498;
wire mux_o_499;
wire mux_o_500;
wire mux_o_501;
wire mux_o_502;
wire mux_o_503;
wire mux_o_504;
wire mux_o_505;
wire mux_o_506;
wire mux_o_507;
wire mux_o_508;
wire mux_o_509;
wire mux_o_510;
wire mux_o_511;
wire mux_o_512;
wire mux_o_513;
wire mux_o_514;
wire mux_o_515;
wire mux_o_516;
wire mux_o_517;
wire mux_o_518;
wire mux_o_519;
wire mux_o_520;
wire mux_o_521;
wire mux_o_522;
wire mux_o_523;
wire mux_o_524;
wire mux_o_525;
wire mux_o_527;
wire mux_o_528;
wire mux_o_529;
wire mux_o_530;
wire mux_o_531;
wire mux_o_532;
wire mux_o_533;
wire mux_o_534;
wire mux_o_535;
wire mux_o_536;
wire mux_o_537;
wire mux_o_538;
wire mux_o_539;
wire mux_o_540;
wire mux_o_541;
wire mux_o_542;
wire mux_o_543;
wire mux_o_544;
wire mux_o_545;
wire mux_o_546;
wire mux_o_547;
wire mux_o_548;
wire mux_o_549;
wire mux_o_550;
wire mux_o_551;
wire mux_o_552;
wire mux_o_553;
wire mux_o_554;
wire mux_o_555;
wire mux_o_556;
wire mux_o_558;
wire mux_o_559;
wire mux_o_560;
wire mux_o_561;
wire mux_o_562;
wire mux_o_563;
wire mux_o_564;
wire mux_o_565;
wire mux_o_566;
wire mux_o_567;
wire mux_o_568;
wire mux_o_569;
wire mux_o_570;
wire mux_o_571;
wire mux_o_572;
wire mux_o_573;
wire mux_o_574;
wire mux_o_575;
wire mux_o_576;
wire mux_o_577;
wire mux_o_578;
wire mux_o_579;
wire mux_o_580;
wire mux_o_581;
wire mux_o_582;
wire mux_o_583;
wire mux_o_584;
wire mux_o_585;
wire mux_o_586;
wire mux_o_587;
wire mux_o_589;
wire mux_o_590;
wire mux_o_591;
wire mux_o_592;
wire mux_o_593;
wire mux_o_594;
wire mux_o_595;
wire mux_o_596;
wire mux_o_597;
wire mux_o_598;
wire mux_o_599;
wire mux_o_600;
wire mux_o_601;
wire mux_o_602;
wire mux_o_603;
wire mux_o_604;
wire mux_o_605;
wire mux_o_606;
wire mux_o_607;
wire mux_o_608;
wire mux_o_609;
wire mux_o_610;
wire mux_o_611;
wire mux_o_612;
wire mux_o_613;
wire mux_o_614;
wire mux_o_615;
wire mux_o_616;
wire mux_o_617;
wire mux_o_618;
wire mux_o_620;
wire mux_o_621;
wire mux_o_622;
wire mux_o_623;
wire mux_o_624;
wire mux_o_625;
wire mux_o_626;
wire mux_o_627;
wire mux_o_628;
wire mux_o_629;
wire mux_o_630;
wire mux_o_631;
wire mux_o_632;
wire mux_o_633;
wire mux_o_634;
wire mux_o_635;
wire mux_o_636;
wire mux_o_637;
wire mux_o_638;
wire mux_o_639;
wire mux_o_640;
wire mux_o_641;
wire mux_o_642;
wire mux_o_643;
wire mux_o_644;
wire mux_o_645;
wire mux_o_646;
wire mux_o_647;
wire mux_o_648;
wire mux_o_649;
wire mux_o_651;
wire mux_o_652;
wire mux_o_653;
wire mux_o_654;
wire mux_o_655;
wire mux_o_656;
wire mux_o_657;
wire mux_o_658;
wire mux_o_659;
wire mux_o_660;
wire mux_o_661;
wire mux_o_662;
wire mux_o_663;
wire mux_o_664;
wire mux_o_665;
wire mux_o_666;
wire mux_o_667;
wire mux_o_668;
wire mux_o_669;
wire mux_o_670;
wire mux_o_671;
wire mux_o_672;
wire mux_o_673;
wire mux_o_674;
wire mux_o_675;
wire mux_o_676;
wire mux_o_677;
wire mux_o_678;
wire mux_o_679;
wire mux_o_680;
wire mux_o_682;
wire mux_o_683;
wire mux_o_684;
wire mux_o_685;
wire mux_o_686;
wire mux_o_687;
wire mux_o_688;
wire mux_o_689;
wire mux_o_690;
wire mux_o_691;
wire mux_o_692;
wire mux_o_693;
wire mux_o_694;
wire mux_o_695;
wire mux_o_696;
wire mux_o_697;
wire mux_o_698;
wire mux_o_699;
wire mux_o_700;
wire mux_o_701;
wire mux_o_702;
wire mux_o_703;
wire mux_o_704;
wire mux_o_705;
wire mux_o_706;
wire mux_o_707;
wire mux_o_708;
wire mux_o_709;
wire mux_o_710;
wire mux_o_711;
wire mux_o_713;
wire mux_o_714;
wire mux_o_715;
wire mux_o_716;
wire mux_o_717;
wire mux_o_718;
wire mux_o_719;
wire mux_o_720;
wire mux_o_721;
wire mux_o_722;
wire mux_o_723;
wire mux_o_724;
wire mux_o_725;
wire mux_o_726;
wire mux_o_727;
wire mux_o_728;
wire mux_o_729;
wire mux_o_730;
wire mux_o_731;
wire mux_o_732;
wire mux_o_733;
wire mux_o_734;
wire mux_o_735;
wire mux_o_736;
wire mux_o_737;
wire mux_o_738;
wire mux_o_739;
wire mux_o_740;
wire mux_o_741;
wire mux_o_742;
wire mux_o_744;
wire mux_o_745;
wire mux_o_746;
wire mux_o_747;
wire mux_o_748;
wire mux_o_749;
wire mux_o_750;
wire mux_o_751;
wire mux_o_752;
wire mux_o_753;
wire mux_o_754;
wire mux_o_755;
wire mux_o_756;
wire mux_o_757;
wire mux_o_758;
wire mux_o_759;
wire mux_o_760;
wire mux_o_761;
wire mux_o_762;
wire mux_o_763;
wire mux_o_764;
wire mux_o_765;
wire mux_o_766;
wire mux_o_767;
wire mux_o_768;
wire mux_o_769;
wire mux_o_770;
wire mux_o_771;
wire mux_o_772;
wire mux_o_773;
wire mux_o_775;
wire mux_o_776;
wire mux_o_777;
wire mux_o_778;
wire mux_o_779;
wire mux_o_780;
wire mux_o_781;
wire mux_o_782;
wire mux_o_783;
wire mux_o_784;
wire mux_o_785;
wire mux_o_786;
wire mux_o_787;
wire mux_o_788;
wire mux_o_789;
wire mux_o_790;
wire mux_o_791;
wire mux_o_792;
wire mux_o_793;
wire mux_o_794;
wire mux_o_795;
wire mux_o_796;
wire mux_o_797;
wire mux_o_798;
wire mux_o_799;
wire mux_o_800;
wire mux_o_801;
wire mux_o_802;
wire mux_o_803;
wire mux_o_804;
wire mux_o_806;
wire mux_o_807;
wire mux_o_808;
wire mux_o_809;
wire mux_o_810;
wire mux_o_811;
wire mux_o_812;
wire mux_o_813;
wire mux_o_814;
wire mux_o_815;
wire mux_o_816;
wire mux_o_817;
wire mux_o_818;
wire mux_o_819;
wire mux_o_820;
wire mux_o_821;
wire mux_o_822;
wire mux_o_823;
wire mux_o_824;
wire mux_o_825;
wire mux_o_826;
wire mux_o_827;
wire mux_o_828;
wire mux_o_829;
wire mux_o_830;
wire mux_o_831;
wire mux_o_832;
wire mux_o_833;
wire mux_o_834;
wire mux_o_835;
wire mux_o_837;
wire mux_o_838;
wire mux_o_839;
wire mux_o_840;
wire mux_o_841;
wire mux_o_842;
wire mux_o_843;
wire mux_o_844;
wire mux_o_845;
wire mux_o_846;
wire mux_o_847;
wire mux_o_848;
wire mux_o_849;
wire mux_o_850;
wire mux_o_851;
wire mux_o_852;
wire mux_o_853;
wire mux_o_854;
wire mux_o_855;
wire mux_o_856;
wire mux_o_857;
wire mux_o_858;
wire mux_o_859;
wire mux_o_860;
wire mux_o_861;
wire mux_o_862;
wire mux_o_863;
wire mux_o_864;
wire mux_o_865;
wire mux_o_866;
wire mux_o_868;
wire mux_o_869;
wire mux_o_870;
wire mux_o_871;
wire mux_o_872;
wire mux_o_873;
wire mux_o_874;
wire mux_o_875;
wire mux_o_876;
wire mux_o_877;
wire mux_o_878;
wire mux_o_879;
wire mux_o_880;
wire mux_o_881;
wire mux_o_882;
wire mux_o_883;
wire mux_o_884;
wire mux_o_885;
wire mux_o_886;
wire mux_o_887;
wire mux_o_888;
wire mux_o_889;
wire mux_o_890;
wire mux_o_891;
wire mux_o_892;
wire mux_o_893;
wire mux_o_894;
wire mux_o_895;
wire mux_o_896;
wire mux_o_897;
wire mux_o_899;
wire mux_o_900;
wire mux_o_901;
wire mux_o_902;
wire mux_o_903;
wire mux_o_904;
wire mux_o_905;
wire mux_o_906;
wire mux_o_907;
wire mux_o_908;
wire mux_o_909;
wire mux_o_910;
wire mux_o_911;
wire mux_o_912;
wire mux_o_913;
wire mux_o_914;
wire mux_o_915;
wire mux_o_916;
wire mux_o_917;
wire mux_o_918;
wire mux_o_919;
wire mux_o_920;
wire mux_o_921;
wire mux_o_922;
wire mux_o_923;
wire mux_o_924;
wire mux_o_925;
wire mux_o_926;
wire mux_o_927;
wire mux_o_928;
wire mux_o_930;
wire mux_o_931;
wire mux_o_932;
wire mux_o_933;
wire mux_o_934;
wire mux_o_935;
wire mux_o_936;
wire mux_o_937;
wire mux_o_938;
wire mux_o_939;
wire mux_o_940;
wire mux_o_941;
wire mux_o_942;
wire mux_o_943;
wire mux_o_944;
wire mux_o_945;
wire mux_o_946;
wire mux_o_947;
wire mux_o_948;
wire mux_o_949;
wire mux_o_950;
wire mux_o_951;
wire mux_o_952;
wire mux_o_953;
wire mux_o_954;
wire mux_o_955;
wire mux_o_956;
wire mux_o_957;
wire mux_o_958;
wire mux_o_959;
wire mux_o_961;
wire mux_o_962;
wire mux_o_963;
wire mux_o_964;
wire mux_o_965;
wire mux_o_966;
wire mux_o_967;
wire mux_o_968;
wire mux_o_969;
wire mux_o_970;
wire mux_o_971;
wire mux_o_972;
wire mux_o_973;
wire mux_o_974;
wire mux_o_975;
wire mux_o_976;
wire mux_o_977;
wire mux_o_978;
wire mux_o_979;
wire mux_o_980;
wire mux_o_981;
wire mux_o_982;
wire mux_o_983;
wire mux_o_984;
wire mux_o_985;
wire mux_o_986;
wire mux_o_987;
wire mux_o_988;
wire mux_o_989;
wire mux_o_990;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT5 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_0.INIT = 32'h00000001;
LUT5 lut_inst_1 (
  .F(lut_f_1),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_1.INIT = 32'h00000002;
LUT5 lut_inst_2 (
  .F(lut_f_2),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_2.INIT = 32'h00000004;
LUT5 lut_inst_3 (
  .F(lut_f_3),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_3.INIT = 32'h00000008;
LUT5 lut_inst_4 (
  .F(lut_f_4),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_4.INIT = 32'h00000010;
LUT5 lut_inst_5 (
  .F(lut_f_5),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_5.INIT = 32'h00000020;
LUT5 lut_inst_6 (
  .F(lut_f_6),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_6.INIT = 32'h00000040;
LUT5 lut_inst_7 (
  .F(lut_f_7),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_7.INIT = 32'h00000080;
LUT5 lut_inst_8 (
  .F(lut_f_8),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_8.INIT = 32'h00000100;
LUT5 lut_inst_9 (
  .F(lut_f_9),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_9.INIT = 32'h00000200;
LUT5 lut_inst_10 (
  .F(lut_f_10),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_10.INIT = 32'h00000400;
LUT5 lut_inst_11 (
  .F(lut_f_11),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_11.INIT = 32'h00000800;
LUT5 lut_inst_12 (
  .F(lut_f_12),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_12.INIT = 32'h00001000;
LUT5 lut_inst_13 (
  .F(lut_f_13),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_13.INIT = 32'h00002000;
LUT5 lut_inst_14 (
  .F(lut_f_14),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_14.INIT = 32'h00004000;
LUT5 lut_inst_15 (
  .F(lut_f_15),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_15.INIT = 32'h00008000;
LUT5 lut_inst_16 (
  .F(lut_f_16),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_16.INIT = 32'h00010000;
LUT5 lut_inst_17 (
  .F(lut_f_17),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_17.INIT = 32'h00020000;
LUT5 lut_inst_18 (
  .F(lut_f_18),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_18.INIT = 32'h00040000;
LUT5 lut_inst_19 (
  .F(lut_f_19),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_19.INIT = 32'h00080000;
LUT5 lut_inst_20 (
  .F(lut_f_20),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_20.INIT = 32'h00100000;
LUT5 lut_inst_21 (
  .F(lut_f_21),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_21.INIT = 32'h00200000;
LUT5 lut_inst_22 (
  .F(lut_f_22),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_22.INIT = 32'h00400000;
LUT5 lut_inst_23 (
  .F(lut_f_23),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_23.INIT = 32'h00800000;
LUT5 lut_inst_24 (
  .F(lut_f_24),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_24.INIT = 32'h01000000;
LUT5 lut_inst_25 (
  .F(lut_f_25),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_25.INIT = 32'h02000000;
LUT5 lut_inst_26 (
  .F(lut_f_26),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_26.INIT = 32'h04000000;
LUT5 lut_inst_27 (
  .F(lut_f_27),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_27.INIT = 32'h08000000;
LUT5 lut_inst_28 (
  .F(lut_f_28),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_28.INIT = 32'h10000000;
LUT5 lut_inst_29 (
  .F(lut_f_29),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_29.INIT = 32'h20000000;
LUT5 lut_inst_30 (
  .F(lut_f_30),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_30.INIT = 32'h40000000;
LUT5 lut_inst_31 (
  .F(lut_f_31),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_31.INIT = 32'h80000000;
SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[15:0],sp_inst_0_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b01;
defparam sp_inst_0.BIT_WIDTH = 16;
defparam sp_inst_0.BLK_SEL = 3'b001;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h000CD1CF358E01EF002F018C002C11AD020F3590020F35F051EF006F2000000D;
defparam sp_inst_0.INIT_RAM_01 = 256'hFD8CE3EC118CFD8C002C102C000C302C002CF9AC118C018011AC01AD000D018C;
defparam sp_inst_0.INIT_RAM_02 = 256'h00000000000000000020800000201800F06300230180200C402C418CA06C442C;
defparam sp_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[15:0],sp_inst_1_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_1}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b01;
defparam sp_inst_1.BIT_WIDTH = 16;
defparam sp_inst_1.BLK_SEL = 3'b001;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'h92A8A2A7B2A6C2A5D2A472B482B392B2A2B1B2B0C2AFD2AEE2ADF2AC0055C435;
defparam sp_inst_1.INIT_RAM_01 = 256'h2DA0818D2DA0418D2DA0218D2DA0118D65A0F18D140C42A352A162AB72AA82A9;
defparam sp_inst_1.INIT_RAM_02 = 256'h140074001C00E0002400C8002C009400340010003C00D0002DA0018D2DA0018D;
defparam sp_inst_1.INIT_RAM_03 = 256'hC2A5D2A472B482B392B2A2B1B2B0C2AFD2AEE2ADF2AC0055040080000DA0018D;
defparam sp_inst_1.INIT_RAM_04 = 256'h0000018C100C40763076C0633800C41542A352A162AB72AA82A992A8A2A7B2A6;
defparam sp_inst_1.INIT_RAM_05 = 256'h102C040C40763076C0630020406330760000042040763076C063002040633076;
defparam sp_inst_1.INIT_RAM_06 = 256'h0000318DB2CC31ADA2CC318DB2CCA2C5B2C48076707680630020406330760000;
defparam sp_inst_1.INIT_RAM_07 = 256'h6076706100008C00D0040185BECCBECC008C8076607670618063002080637076;
defparam sp_inst_1.INIT_RAM_08 = 256'h300C72CC1D8072CC258042CC42C752C662C572C4C076A076B061406300208063;
defparam sp_inst_1.INIT_RAM_09 = 256'hC2CEB2CD5DCC00070980B1AE92CD52CC5000B2C092CC72CC0C0087FFB40492CC;
defparam sp_inst_1.INIT_RAM_0A = 256'hB2CEB2CD62CCB19F92CCB2CC058CB2CC92CC000709A035CC92CE52CDC1AC35CD;
defparam sp_inst_1.INIT_RAM_0B = 256'h000C0800C18C31ACC2CDFD8CA2CC1D8DB2CCA2CD7400A2CC31CC358CB5CE31AD;
defparam sp_inst_1.INIT_RAM_0C = 256'hA2CC97FF0184818C5D8C818C82CC1400818CC18C818C82CC198D240C82CD82CC;
defparam sp_inst_1.INIT_RAM_0D = 256'h300072C4C076A076B06140630020C063A076B0610184000C8C0CA2CCA2CCFD8C;
defparam sp_inst_1.INIT_RAM_0E = 256'hC59FBECCBECC018C72CC72CC058C72CC33FF0184BECC3FFF34040DAC280CBECD;
defparam sp_inst_1.INIT_RAM_0F = 256'h52C942C832C722C612C532C40076E076F06180630020C063A076B0610184000C;
defparam sp_inst_1.INIT_RAM_10 = 256'h940C8ECD8ECC018C31AC32CDB2CC3000B2C0A2CC72CC72CC918C82CC72CB62CA;
defparam sp_inst_1.INIT_RAM_11 = 256'h018C31ACD18C002C898DADAC4C0D6D8C018C31AC32CD058CB2CC92CC040CE5AC;
defparam sp_inst_1.INIT_RAM_12 = 256'h0184818C018CA2CC9800B2CC058CB2CCA2CC118CA2CCDBFF0184018CA2CC0180;
defparam sp_inst_1.INIT_RAM_13 = 256'hA2CC13FF018492C528060007018CA2CC6800B2CC058CB2CCA2CC118CA2CC0FFF;
defparam sp_inst_1.INIT_RAM_14 = 256'hA2CC118CA2CCDBFF018492C528060407018CA2CC3000B2CC058CB2CCA2CC118C;
defparam sp_inst_1.INIT_RAM_15 = 256'h058CB2CCA2CC118CA2CCA3FF018492C520060007018CA2CCF800B2CC058CB2CC;
defparam sp_inst_1.INIT_RAM_16 = 256'h8800B2CC058CB2CCA2CC118CA2CC6BFF018492C508060007018CA2CCC000B2CC;
defparam sp_inst_1.INIT_RAM_17 = 256'hD3FF94045000B2CC058CB2CCA2CC118CA2CC33FF018492C540060007018CA2CC;
defparam sp_inst_1.INIT_RAM_18 = 256'h31CC32CE058CB2CC31AD280C92CD3C0092C0B2CC058CB2CC3800B2CC058CB2CC;
defparam sp_inst_1.INIT_RAM_19 = 256'h058CB2CCD98DC00C018D31AC32CD058CB2CCB2CC058CB2CC92CC31AC418C018C;
defparam sp_inst_1.INIT_RAM_1A = 256'h018C31CC32CE058CB2CC31AD280C92CD3C0092C0BBFF958DE40C018D31AC32CD;
defparam sp_inst_1.INIT_RAM_1B = 256'h32CD058CB2CC5D8DC00C018D31AC32CD058CB2CCB2CC058CB2CC92CC31AC418C;
defparam sp_inst_1.INIT_RAM_1C = 256'h01848ECC9BFF34040DAC280C8ECD24000000B7FF94043FFF958DE40C018D31AC;
defparam sp_inst_1.INIT_RAM_1D = 256'h806300208063E076F0610184000CC59F018C31AC32CDB2CCB2CC058CB2CC8FFF;
defparam sp_inst_1.INIT_RAM_1E = 256'h70760000018DAECDB2CCF19F818C818C158CB2CC0000AECC00ACB2C480767076;
defparam sp_inst_1.INIT_RAM_1F = 256'hC076B07640630020406330760000D18DA9ADB4ADD60C40763076C06300208063;
defparam sp_inst_1.INIT_RAM_20 = 256'h018E300C31CCB2CC040E018DD60C318062CCB2CC72CC698D7C0C72CD62C572C4;
defparam sp_inst_1.INIT_RAM_21 = 256'h818C72CC6800018D39ADD60C018E31CCB2CC040E018DD60C9000018DB9ADD60C;
defparam sp_inst_1.INIT_RAM_22 = 256'h418DD60C2800418DB9ADD60C018E300C31CCB2CC040E418DD60C318062CCB2CC;
defparam sp_inst_1.INIT_RAM_23 = 256'h62C572C4C076B07640630020C063B0760000418D39ADD60C018E31CCB2CC040E;
defparam sp_inst_1.INIT_RAM_24 = 256'hB9ADD60C018E300C31CCB2CC040E118DD60C318062CCB2CC72CC698D7C0C72CD;
defparam sp_inst_1.INIT_RAM_25 = 256'h62CCB2CC818C72CC6800118D39ADD60C018E31CCB2CC040E118DD60C9000118D;
defparam sp_inst_1.INIT_RAM_26 = 256'hB2CC040E518DD60C2800518DB9ADD60C018E300C31CCB2CC040E518DD60C3180;
defparam sp_inst_1.INIT_RAM_27 = 256'h018DDA0CB2C072C4C076B07640630020C063B0760000518D39ADD60C018E31CC;
defparam sp_inst_1.INIT_RAM_28 = 256'hB2C48076707680630020C063B0760184B2CCB2C00800B2CC040C1180B1AC72CC;
defparam sp_inst_1.INIT_RAM_29 = 256'h0000018D81AD05AD0D8CD40C818D018C0D8CD40C018D35CDB2CDDA0C018EDA0C;
defparam sp_inst_1.INIT_RAM_2A = 256'hFFC40185BECC018D040D718CFFCCBECC008C8076607670618063002080637076;
defparam sp_inst_1.INIT_RAM_2B = 256'hB2CD018CB2CCAECC00ACB2C48076707680630020806360767061000018002084;
defparam sp_inst_1.INIT_RAM_2C = 256'h3180B2CC0DAC118CB2CC318DB2CC318DB2CC058D318CB2CC018DAECD358C31AD;
defparam sp_inst_1.INIT_RAM_2D = 256'h218CB2CC418DB2CC118DB2CC458D118CB2CC418DB2CC418DB2CC058D418CB2CC;
defparam sp_inst_1.INIT_RAM_2E = 256'h7061806300208063707600002180B2CC0DAC118CB2CC218DB2CC218DB2CC058D;
defparam sp_inst_1.INIT_RAM_2F = 256'h0405FFFF4C0404050BFF4804040517FF3404040523FF0404040563FF80766076;
defparam sp_inst_1.INIT_RAM_30 = 256'h98040405C3FF94040405CFFF90040405DBFF8C040405E7FF88040405F3FF5004;
defparam sp_inst_1.INIT_RAM_31 = 256'hB2CC00000000000000001400B2CC918C1C6C9FFFA0040405ABFF9C040405B7FF;
defparam sp_inst_1.INIT_RAM_32 = 256'h040537FF4C04040543FF480404054FFF340404055BFF04040405E59FB2CDFD8D;
defparam sp_inst_1.INIT_RAM_33 = 256'h98040405FBFF9404040507FF9004040513FF8C0404051FFF880404052BFF5004;
defparam sp_inst_1.INIT_RAM_34 = 256'hA2CC00000000000000001400A2CC918C1C6CD7FFA0040405E3FF9C040405EFFF;
defparam sp_inst_1.INIT_RAM_35 = 256'h000577FF4C04000583FF480400058FFF340400059BFF04040005E59FA2CDFD8D;
defparam sp_inst_1.INIT_RAM_36 = 256'h980400053BFF9404000547FF9004000553FF8C0400055FFF880400056BFF5004;
defparam sp_inst_1.INIT_RAM_37 = 256'h92CC0000000000000000140092CC918C1C6C17FFA004000523FF9C0400052FFF;
defparam sp_inst_1.INIT_RAM_38 = 256'hD60C0405A7FF208400244C05A0C60026407620763061C06383FFE59F92CDFD8D;
defparam sp_inst_1.INIT_RAM_39 = 256'hF08400246005D0C60026407620763061C063002040632076306100004FFF8184;
defparam sp_inst_1.INIT_RAM_3A = 256'h00C60026407620763061C0630020406320763061000003FF8184D60C08055BFF;
defparam sp_inst_1.INIT_RAM_3B = 256'h20763061C06300204063207630610000B7FF8184D60C10050FFFC08400247405;
defparam sp_inst_1.INIT_RAM_3C = 256'h002040632076306100006BFF8184D60C2005C3FF90840024880530C600264076;
defparam sp_inst_1.INIT_RAM_3D = 256'h306100001FFF8184D60C400577FF608400249C0560C60026407620763061C063;
defparam sp_inst_1.INIT_RAM_3E = 256'h8184D60C80052BFF30840024B00590C60026407620763061C063002040632076;
defparam sp_inst_1.INIT_RAM_3F = 256'hDFFF00840024C405C0C60026407620763061C06300204063207630610000D3FF;

SP sp_inst_2 (
    .DO({sp_inst_2_dout_w[15:0],sp_inst_2_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_2}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_2.READ_MODE = 1'b0;
defparam sp_inst_2.WRITE_MODE = 2'b01;
defparam sp_inst_2.BIT_WIDTH = 16;
defparam sp_inst_2.BLK_SEL = 3'b001;
defparam sp_inst_2.RESET_MODE = "SYNC";
defparam sp_inst_2.INIT_RAM_00 = 256'hDC05F0C60026407620763061C0630020406320763061000087FF8184D60C0005;
defparam sp_inst_2.INIT_RAM_01 = 256'h407620763061C063002040632076306100003BFF8184D60C000593FFD0840024;
defparam sp_inst_2.INIT_RAM_02 = 256'hC06300204063207630610000EFFF8184D60C000547FFA0840024F00520C60026;
defparam sp_inst_2.INIT_RAM_03 = 256'h207630610000A3FF8184D60C0005FBFF70840024080550C60026407620763061;
defparam sp_inst_2.INIT_RAM_04 = 256'h57FF8184D60C0005AFFF40840024200580C60026407620763061C06300204063;
defparam sp_inst_2.INIT_RAM_05 = 256'h000563FF108400243805B0C60026407620763061C06300204063207630610000;
defparam sp_inst_2.INIT_RAM_06 = 256'h00244C05E0C60026407620763061C063002040632076306100000BFF8184D60C;
defparam sp_inst_2.INIT_RAM_07 = 256'h0026407620763061C06300204063207630610000BFFF8184D60C002517FFE084;
defparam sp_inst_2.INIT_RAM_08 = 256'h3061C0630020406320763061000073FF8184D60C0045CBFFB0840024600510C6;
defparam sp_inst_2.INIT_RAM_09 = 256'h406320763061000027FF8184D60C00857FFF80840024780540C6002640762076;
defparam sp_inst_2.INIT_RAM_0A = 256'h0000DBFF8184D60C010533FF50840024900570C60026407620763061C0630020;
defparam sp_inst_2.INIT_RAM_0B = 256'hD60C0205E7FF20840024AC05A0C60026407620763061C0630020406320763061;
defparam sp_inst_2.INIT_RAM_0C = 256'hF0840024C405D0C60026407620763061C063002040632076306100008FFF8184;
defparam sp_inst_2.INIT_RAM_0D = 256'h00C60026407620763061C0630020406320763061000043FF8184D60C04059BFF;
defparam sp_inst_2.INIT_RAM_0E = 256'h20763061C06300204063207630610000F7FF8184D60C08054FFFC0840024DC05;
defparam sp_inst_2.INIT_RAM_0F = 256'h00204063207630610000ABFF8184D60C100503FF90840024F40530C600264076;
defparam sp_inst_2.INIT_RAM_10 = 256'h306100005FFF8184D60C2005B7FF608400240C0560C60026407620763061C063;
defparam sp_inst_2.INIT_RAM_11 = 256'h8184D60C40056BFF30840024200590C60026407620763061C063002040632076;
defparam sp_inst_2.INIT_RAM_12 = 256'h1FFF008400243405C0C60026407620763061C0630020406320763061000013FF;
defparam sp_inst_2.INIT_RAM_13 = 256'h4C05F0C60026407620763061C06300204063207630610000C7FF8184D60C8005;
defparam sp_inst_2.INIT_RAM_14 = 256'h407620763061C063002040632076306100007BFF8184D60C0005D3FFD0840004;
defparam sp_inst_2.INIT_RAM_15 = 256'hC063002040632076306100002FFF8184D60C000587FFA0840004640520C60026;
defparam sp_inst_2.INIT_RAM_16 = 256'h207630610000E3FF8184D60C00053BFF708400047C0550C60026407620763061;
defparam sp_inst_2.INIT_RAM_17 = 256'h97FF8184D60C0005EFFF40840004940580C60026407620763061C06300204063;
defparam sp_inst_2.INIT_RAM_18 = 256'h0005A3FF10840004AC05B0C60026407620763061C06300204063207630610000;
defparam sp_inst_2.INIT_RAM_19 = 256'h0004C405E0C60026407620763061C063002040632076306100004BFF8184D60C;
defparam sp_inst_2.INIT_RAM_1A = 256'h0026407620763061C06300204063207630610000FFFF8184D60C000557FFE084;
defparam sp_inst_2.INIT_RAM_1B = 256'h3061C06300204063207630610000B3FF8184D60C00050BFFB0840004E00510C6;
defparam sp_inst_2.INIT_RAM_1C = 256'h406320763061000067FF8184D60C0005BFFF80840004F80540C6002640762076;
defparam sp_inst_2.INIT_RAM_1D = 256'h00001BFF8184D60C000573FF50840004100570C60026407620763061C0630020;
defparam sp_inst_2.INIT_RAM_1E = 256'h0004C00560C60026018D000DF18CD60C80766076706180630020406320763061;
defparam sp_inst_2.INIT_RAM_1F = 256'hB2C00000A2CCB1AC92CCA2CD92CC018C818CD60CA2CC318C818CD60C17FFE084;
defparam sp_inst_2.INIT_RAM_20 = 256'hB2CC058CB2CC0181018C31AC898CB2CCB1AD000D2180058CB1ACB2CCA2CD4000;
defparam sp_inst_2.INIT_RAM_21 = 256'h018D020DF18CD60C807660767061806300208063607670610000BD8D7C0CB2CD;
defparam sp_inst_2.INIT_RAM_22 = 256'h118CD68C8076607670618063002080636076706100003BFFB2CC018C118CD60C;
defparam sp_inst_2.INIT_RAM_23 = 256'hD68C018D040DF18CD60CB6CC3D8C818C018C118CD68CBACCFD8C818CC18C018C;
defparam sp_inst_2.INIT_RAM_24 = 256'h80767076806300208063607670610000BFFFA08400040185BACC018D3C0D118C;
defparam sp_inst_2.INIT_RAM_25 = 256'h80766076706180630020806370760000BECC018C098CD18C018D080DF18CD60C;
defparam sp_inst_2.INIT_RAM_26 = 256'h400CB2CD018DB5CDF00DF18CD60C018E118CD60CB2CC7D8CCD8C018C118CD60C;
defparam sp_inst_2.INIT_RAM_27 = 256'h00043C000180118CD60CF3FFF08400040180018C31ACE18C000C898DB2CC718D;
defparam sp_inst_2.INIT_RAM_28 = 256'h60767061000000000800018DB5CDFDADFEED118CD60C018E118CD60CD7FF2084;
defparam sp_inst_2.INIT_RAM_29 = 256'h008C6FFF00042980058CBECCBECC018C158CD40C807660767061806300208063;
defparam sp_inst_2.INIT_RAM_2A = 256'h608400040185BACCBACC018CD10C3580118CBECC47FF70840004ABFF00041980;
defparam sp_inst_2.INIT_RAM_2B = 256'h0D8CD40C9BFF0184B6CCB6CC018CD00C2D80218CBECC018D100D0D8CD40C1BFF;
defparam sp_inst_2.INIT_RAM_2C = 256'h33FF407620763061C06300208063607670610000018DFC0D0D8CD40C018D200D;
defparam sp_inst_2.INIT_RAM_2D = 256'h17141714171417141714171415F80020406320763061000003FF93FF90840004;
defparam sp_inst_2.INIT_RAM_2E = 256'h1714171416981698169816981698169816981698169816101714171417141714;
defparam sp_inst_2.INIT_RAM_2F = 256'h1714171417141714171417141714171417141714171417141714171417141714;
defparam sp_inst_2.INIT_RAM_30 = 256'h1714171417141714171417141714171417141714171417141714171417141714;
defparam sp_inst_2.INIT_RAM_31 = 256'h1714171417141714171417141714151814B01588171417141714171417141714;
defparam sp_inst_2.INIT_RAM_32 = 256'h656E20200A0D15C01714171414E0171414841714171415C01550171417141714;
defparam sp_inst_2.INIT_RAM_33 = 256'h2D0A0D0A2E2E2E2E2E2E544E54462E2E2E2E2E2E2E0A00003E2073256E756425;
defparam sp_inst_2.INIT_RAM_34 = 256'h2E2E2E2E2E2E4C495F542E2E2E2E2E2E2E0A000A7830656E68434B3A49686F74;
defparam sp_inst_2.INIT_RAM_35 = 256'h6165207269546C6168706550000D2E2E2E2E2E2E2E432E2E2E2E2E2E2E0A0D0A;
defparam sp_inst_2.INIT_RAM_36 = 256'h747072656920656C726554206F430000257876632031617500002E7472726E69;
defparam sp_inst_2.INIT_RAM_37 = 256'h223821EC21A02154210820BC207020241FD81F8C1F401EF41EA81E5C1E10000A;
defparam sp_inst_2.INIT_RAM_38 = 256'h26F826AC2660261425C8257C253024E42498244C240023B42368231C22D02284;
defparam sp_inst_2.INIT_RAM_39 = 256'h2A302A302A302A302A302A302A302A302A302A302A302A302A3029E02A302744;
defparam sp_inst_2.INIT_RAM_3A = 256'h675F7865656C61687269616F675F7865656C61687269616F675F786529FC2A30;
defparam sp_inst_2.INIT_RAM_3B = 256'h656C61687269616F675F7865656C61687269616F675F7865656C61687269616F;
defparam sp_inst_2.INIT_RAM_3C = 256'h7269616F675F7865656C61687269616F675F7865656C61687269616F675F7865;
defparam sp_inst_2.INIT_RAM_3D = 256'h675F7865656C61687269626F675F7865656C61687269626F675F7865656C6168;
defparam sp_inst_2.INIT_RAM_3E = 256'h656C61687269626F675F7865656C61687269626F675F7865656C61687269626F;
defparam sp_inst_2.INIT_RAM_3F = 256'h7269626F675F7865656C61687269626F675F7865656C61687269626F675F7865;

SP sp_inst_3 (
    .DO({sp_inst_3_dout_w[15:0],sp_inst_3_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_3}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_3.READ_MODE = 1'b0;
defparam sp_inst_3.WRITE_MODE = 2'b01;
defparam sp_inst_3.BIT_WIDTH = 16;
defparam sp_inst_3.BLK_SEL = 3'b001;
defparam sp_inst_3.RESET_MODE = "SYNC";
defparam sp_inst_3.INIT_RAM_00 = 256'h675F7865656C61687269636F675F7865656C61687269636F675F7865656C6168;
defparam sp_inst_3.INIT_RAM_01 = 256'h656C61687269636F675F7865656C61687269636F675F7865656C61687269636F;
defparam sp_inst_3.INIT_RAM_02 = 256'h7269636F675F7865656C61687269636F675F7865656C61687269636F675F7865;
defparam sp_inst_3.INIT_RAM_03 = 256'h675F7865656C61687269646F675F7865656C61687269646F675F7865656C6168;
defparam sp_inst_3.INIT_RAM_04 = 256'h656C61687269646F675F7865656C61687269646F675F7865656C61687269646F;
defparam sp_inst_3.INIT_RAM_05 = 256'h7269646F675F7865656C61687269646F675F7865656C61687269646F675F7865;
defparam sp_inst_3.INIT_RAM_06 = 256'h00000000000000000000000000000000000000000000656C61687865656C6168;
defparam sp_inst_3.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_4 (
    .DO({sp_inst_4_dout_w[15:0],sp_inst_4_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_4}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_4.READ_MODE = 1'b0;
defparam sp_inst_4.WRITE_MODE = 2'b01;
defparam sp_inst_4.BIT_WIDTH = 16;
defparam sp_inst_4.BLK_SEL = 3'b001;
defparam sp_inst_4.RESET_MODE = "SYNC";
defparam sp_inst_4.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_4.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_5 (
    .DO({sp_inst_5_dout_w[15:0],sp_inst_5_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_5}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_5.READ_MODE = 1'b0;
defparam sp_inst_5.WRITE_MODE = 2'b01;
defparam sp_inst_5.BIT_WIDTH = 16;
defparam sp_inst_5.BLK_SEL = 3'b001;
defparam sp_inst_5.RESET_MODE = "SYNC";
defparam sp_inst_5.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_6 (
    .DO({sp_inst_6_dout_w[15:0],sp_inst_6_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_6}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_6.READ_MODE = 1'b0;
defparam sp_inst_6.WRITE_MODE = 2'b01;
defparam sp_inst_6.BIT_WIDTH = 16;
defparam sp_inst_6.BLK_SEL = 3'b001;
defparam sp_inst_6.RESET_MODE = "SYNC";
defparam sp_inst_6.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_7 (
    .DO({sp_inst_7_dout_w[15:0],sp_inst_7_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_7}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_7.READ_MODE = 1'b0;
defparam sp_inst_7.WRITE_MODE = 2'b01;
defparam sp_inst_7.BIT_WIDTH = 16;
defparam sp_inst_7.BLK_SEL = 3'b001;
defparam sp_inst_7.RESET_MODE = "SYNC";
defparam sp_inst_7.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_8 (
    .DO({sp_inst_8_dout_w[15:0],sp_inst_8_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_8}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_8.READ_MODE = 1'b0;
defparam sp_inst_8.WRITE_MODE = 2'b01;
defparam sp_inst_8.BIT_WIDTH = 16;
defparam sp_inst_8.BLK_SEL = 3'b001;
defparam sp_inst_8.RESET_MODE = "SYNC";
defparam sp_inst_8.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_9 (
    .DO({sp_inst_9_dout_w[15:0],sp_inst_9_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_9}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_9.READ_MODE = 1'b0;
defparam sp_inst_9.WRITE_MODE = 2'b01;
defparam sp_inst_9.BIT_WIDTH = 16;
defparam sp_inst_9.BLK_SEL = 3'b001;
defparam sp_inst_9.RESET_MODE = "SYNC";
defparam sp_inst_9.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_9.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_10 (
    .DO({sp_inst_10_dout_w[15:0],sp_inst_10_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_10}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_10.READ_MODE = 1'b0;
defparam sp_inst_10.WRITE_MODE = 2'b01;
defparam sp_inst_10.BIT_WIDTH = 16;
defparam sp_inst_10.BLK_SEL = 3'b001;
defparam sp_inst_10.RESET_MODE = "SYNC";
defparam sp_inst_10.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_10.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_11 (
    .DO({sp_inst_11_dout_w[15:0],sp_inst_11_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_11}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_11.READ_MODE = 1'b0;
defparam sp_inst_11.WRITE_MODE = 2'b01;
defparam sp_inst_11.BIT_WIDTH = 16;
defparam sp_inst_11.BLK_SEL = 3'b001;
defparam sp_inst_11.RESET_MODE = "SYNC";
defparam sp_inst_11.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_12 (
    .DO({sp_inst_12_dout_w[15:0],sp_inst_12_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_12}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_12.READ_MODE = 1'b0;
defparam sp_inst_12.WRITE_MODE = 2'b01;
defparam sp_inst_12.BIT_WIDTH = 16;
defparam sp_inst_12.BLK_SEL = 3'b001;
defparam sp_inst_12.RESET_MODE = "SYNC";
defparam sp_inst_12.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_12.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_13 (
    .DO({sp_inst_13_dout_w[15:0],sp_inst_13_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_13}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_13.READ_MODE = 1'b0;
defparam sp_inst_13.WRITE_MODE = 2'b01;
defparam sp_inst_13.BIT_WIDTH = 16;
defparam sp_inst_13.BLK_SEL = 3'b001;
defparam sp_inst_13.RESET_MODE = "SYNC";
defparam sp_inst_13.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_13.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_14 (
    .DO({sp_inst_14_dout_w[15:0],sp_inst_14_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_14}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_14.READ_MODE = 1'b0;
defparam sp_inst_14.WRITE_MODE = 2'b01;
defparam sp_inst_14.BIT_WIDTH = 16;
defparam sp_inst_14.BLK_SEL = 3'b001;
defparam sp_inst_14.RESET_MODE = "SYNC";
defparam sp_inst_14.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_14.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_15 (
    .DO({sp_inst_15_dout_w[15:0],sp_inst_15_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_15}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_15.READ_MODE = 1'b0;
defparam sp_inst_15.WRITE_MODE = 2'b01;
defparam sp_inst_15.BIT_WIDTH = 16;
defparam sp_inst_15.BLK_SEL = 3'b001;
defparam sp_inst_15.RESET_MODE = "SYNC";
defparam sp_inst_15.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_15.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_16 (
    .DO({sp_inst_16_dout_w[15:0],sp_inst_16_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_16}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_16.READ_MODE = 1'b0;
defparam sp_inst_16.WRITE_MODE = 2'b01;
defparam sp_inst_16.BIT_WIDTH = 16;
defparam sp_inst_16.BLK_SEL = 3'b001;
defparam sp_inst_16.RESET_MODE = "SYNC";
defparam sp_inst_16.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_17 (
    .DO({sp_inst_17_dout_w[15:0],sp_inst_17_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_17}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_17.READ_MODE = 1'b0;
defparam sp_inst_17.WRITE_MODE = 2'b01;
defparam sp_inst_17.BIT_WIDTH = 16;
defparam sp_inst_17.BLK_SEL = 3'b001;
defparam sp_inst_17.RESET_MODE = "SYNC";
defparam sp_inst_17.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_17.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_18 (
    .DO({sp_inst_18_dout_w[15:0],sp_inst_18_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_18}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_18.READ_MODE = 1'b0;
defparam sp_inst_18.WRITE_MODE = 2'b01;
defparam sp_inst_18.BIT_WIDTH = 16;
defparam sp_inst_18.BLK_SEL = 3'b001;
defparam sp_inst_18.RESET_MODE = "SYNC";
defparam sp_inst_18.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_18.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_19 (
    .DO({sp_inst_19_dout_w[15:0],sp_inst_19_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_19}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_19.READ_MODE = 1'b0;
defparam sp_inst_19.WRITE_MODE = 2'b01;
defparam sp_inst_19.BIT_WIDTH = 16;
defparam sp_inst_19.BLK_SEL = 3'b001;
defparam sp_inst_19.RESET_MODE = "SYNC";
defparam sp_inst_19.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_19.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_20 (
    .DO({sp_inst_20_dout_w[15:0],sp_inst_20_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_20}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_20.READ_MODE = 1'b0;
defparam sp_inst_20.WRITE_MODE = 2'b01;
defparam sp_inst_20.BIT_WIDTH = 16;
defparam sp_inst_20.BLK_SEL = 3'b001;
defparam sp_inst_20.RESET_MODE = "SYNC";
defparam sp_inst_20.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_20.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_21 (
    .DO({sp_inst_21_dout_w[15:0],sp_inst_21_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_21}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_21.READ_MODE = 1'b0;
defparam sp_inst_21.WRITE_MODE = 2'b01;
defparam sp_inst_21.BIT_WIDTH = 16;
defparam sp_inst_21.BLK_SEL = 3'b001;
defparam sp_inst_21.RESET_MODE = "SYNC";
defparam sp_inst_21.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_21.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_22 (
    .DO({sp_inst_22_dout_w[15:0],sp_inst_22_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_22}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_22.READ_MODE = 1'b0;
defparam sp_inst_22.WRITE_MODE = 2'b01;
defparam sp_inst_22.BIT_WIDTH = 16;
defparam sp_inst_22.BLK_SEL = 3'b001;
defparam sp_inst_22.RESET_MODE = "SYNC";
defparam sp_inst_22.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_23 (
    .DO({sp_inst_23_dout_w[15:0],sp_inst_23_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_23}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_23.READ_MODE = 1'b0;
defparam sp_inst_23.WRITE_MODE = 2'b01;
defparam sp_inst_23.BIT_WIDTH = 16;
defparam sp_inst_23.BLK_SEL = 3'b001;
defparam sp_inst_23.RESET_MODE = "SYNC";
defparam sp_inst_23.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_23.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_24 (
    .DO({sp_inst_24_dout_w[15:0],sp_inst_24_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_24}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_24.READ_MODE = 1'b0;
defparam sp_inst_24.WRITE_MODE = 2'b01;
defparam sp_inst_24.BIT_WIDTH = 16;
defparam sp_inst_24.BLK_SEL = 3'b001;
defparam sp_inst_24.RESET_MODE = "SYNC";
defparam sp_inst_24.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_25 (
    .DO({sp_inst_25_dout_w[15:0],sp_inst_25_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_25}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_25.READ_MODE = 1'b0;
defparam sp_inst_25.WRITE_MODE = 2'b01;
defparam sp_inst_25.BIT_WIDTH = 16;
defparam sp_inst_25.BLK_SEL = 3'b001;
defparam sp_inst_25.RESET_MODE = "SYNC";
defparam sp_inst_25.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_25.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_26 (
    .DO({sp_inst_26_dout_w[15:0],sp_inst_26_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_26}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_26.READ_MODE = 1'b0;
defparam sp_inst_26.WRITE_MODE = 2'b01;
defparam sp_inst_26.BIT_WIDTH = 16;
defparam sp_inst_26.BLK_SEL = 3'b001;
defparam sp_inst_26.RESET_MODE = "SYNC";
defparam sp_inst_26.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_26.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_27 (
    .DO({sp_inst_27_dout_w[15:0],sp_inst_27_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_27}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_27.READ_MODE = 1'b0;
defparam sp_inst_27.WRITE_MODE = 2'b01;
defparam sp_inst_27.BIT_WIDTH = 16;
defparam sp_inst_27.BLK_SEL = 3'b001;
defparam sp_inst_27.RESET_MODE = "SYNC";
defparam sp_inst_27.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_27.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_28 (
    .DO({sp_inst_28_dout_w[15:0],sp_inst_28_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_28}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_28.READ_MODE = 1'b0;
defparam sp_inst_28.WRITE_MODE = 2'b01;
defparam sp_inst_28.BIT_WIDTH = 16;
defparam sp_inst_28.BLK_SEL = 3'b001;
defparam sp_inst_28.RESET_MODE = "SYNC";
defparam sp_inst_28.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_28.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_29 (
    .DO({sp_inst_29_dout_w[15:0],sp_inst_29_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_29}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_29.READ_MODE = 1'b0;
defparam sp_inst_29.WRITE_MODE = 2'b01;
defparam sp_inst_29.BIT_WIDTH = 16;
defparam sp_inst_29.BLK_SEL = 3'b001;
defparam sp_inst_29.RESET_MODE = "SYNC";
defparam sp_inst_29.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_29.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_30 (
    .DO({sp_inst_30_dout_w[15:0],sp_inst_30_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_30}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_30.READ_MODE = 1'b0;
defparam sp_inst_30.WRITE_MODE = 2'b01;
defparam sp_inst_30.BIT_WIDTH = 16;
defparam sp_inst_30.BLK_SEL = 3'b001;
defparam sp_inst_30.RESET_MODE = "SYNC";
defparam sp_inst_30.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_30.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_31 (
    .DO({sp_inst_31_dout_w[15:0],sp_inst_31_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_31}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_31.READ_MODE = 1'b0;
defparam sp_inst_31.WRITE_MODE = 2'b01;
defparam sp_inst_31.BIT_WIDTH = 16;
defparam sp_inst_31.BLK_SEL = 3'b001;
defparam sp_inst_31.RESET_MODE = "SYNC";
defparam sp_inst_31.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_31.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_32 (
    .DO({sp_inst_32_dout_w[15:0],sp_inst_32_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_32.READ_MODE = 1'b0;
defparam sp_inst_32.WRITE_MODE = 2'b01;
defparam sp_inst_32.BIT_WIDTH = 16;
defparam sp_inst_32.BLK_SEL = 3'b001;
defparam sp_inst_32.RESET_MODE = "SYNC";
defparam sp_inst_32.INIT_RAM_00 = 256'h15005FFF00100380150003801500028029800010288000100386143850000015;
defparam sp_inst_32.INIT_RAM_01 = 256'h03BF15FF040003BF140004000015040014385FFF028029805800038015000380;
defparam sp_inst_32.INIT_RAM_02 = 256'h00000000000000004C0006484C00541B03BD1500040003800406038814EC0406;
defparam sp_inst_32.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_32.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_33 (
    .DO({sp_inst_33_dout_w[15:0],sp_inst_33_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_1}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_33.READ_MODE = 1'b0;
defparam sp_inst_33.WRITE_MODE = 2'b01;
defparam sp_inst_33.BIT_WIDTH = 16;
defparam sp_inst_33.BLK_SEL = 3'b001;
defparam sp_inst_33.RESET_MODE = "SYNC";
defparam sp_inst_33.INIT_RAM_00 = 256'h29BE29BE29BE29BE29BE29BF29BF29BF29BF29BF29BF29BF29BF29BF15000400;
defparam sp_inst_33.INIT_RAM_01 = 256'h440003404400034044000340440003404000036E040029BE29BE29BE29BE29BE;
defparam sp_inst_33.INIT_RAM_02 = 256'h5000541A50005416500054185000541850005418500054174400036044000342;
defparam sp_inst_33.INIT_RAM_03 = 256'h28BE28BE28BF28BF28BF28BF28BF28BF28BF28BF28BF15005000541940000341;
defparam sp_inst_33.INIT_RAM_04 = 256'h0340040003800280298002BF0648040028BE28BE28BE28BE28BE28BE28BE28BE;
defparam sp_inst_33.INIT_RAM_05 = 256'h040103800280298002BF4C0002802880034004010280298002BF4C0002802880;
defparam sp_inst_33.INIT_RAM_06 = 256'h0340298028BF001528BF288028BF29BF29BF0280298002BF4C00028028800340;
defparam sp_inst_33.INIT_RAM_07 = 256'h2880288003405405157F00152A3F293F001502802980298002BF4C0002802880;
defparam sp_inst_33.INIT_RAM_08 = 256'h001128BE640028BE400028BE29BE29BE29BE29BE02812981298102BE4C000280;
defparam sp_inst_33.INIT_RAM_09 = 256'h02BF28BF0000002A5C00002128BF28BE500029BF29BF28BE500057FF028029BF;
defparam sp_inst_33.INIT_RAM_0A = 256'h28BF28BF28BE47FF28BF29BF028028BF29BF002A5C00002128BF28BE293E0010;
defparam sp_inst_33.INIT_RAM_0B = 256'h00155000283E001002BF02BF28BF600028BF28BF500029BF0015001300130012;
defparam sp_inst_33.INIT_RAM_0C = 256'h28BF57FE001500670281006728BF500000670280006728BF6000028028BF29BF;
defparam sp_inst_33.INIT_RAM_0D = 256'h500029BF02802980298002BF4C000281288128810015001563FF28BF29BF02BF;
defparam sp_inst_33.INIT_RAM_0E = 256'h47FF283F293F2A0028BF29BF028028BF57FE00152A3F57FE02805C000280283F;
defparam sp_inst_33.INIT_RAM_0F = 256'h2980298029802980298029BF02812980298002BE4C0002802880288000150015;
defparam sp_inst_33.INIT_RAM_10 = 256'h0280283F293F2A00001028BF28BF500329BF29BF28BF29BF02BF028029802980;
defparam sp_inst_33.INIT_RAM_11 = 256'h28800010029B1C0000406802028102BF2800001028BF028028BF29BF02805C02;
defparam sp_inst_33.INIT_RAM_12 = 256'h00150067288028BF500229BF028028BF29BF028028BF57FE0015288028BF4C00;
defparam sp_inst_33.INIT_RAM_13 = 256'h28BF57FD001528BF02800015288028BF500229BF028028BF29BF028028BF57FD;
defparam sp_inst_33.INIT_RAM_14 = 256'h29BF028028BF57FC001528BF02800280288028BF500229BF028028BF29BF0280;
defparam sp_inst_33.INIT_RAM_15 = 256'h028028BF29BF028028BF57FC001528BF02800015288028BF500129BF028028BF;
defparam sp_inst_33.INIT_RAM_16 = 256'h500129BF028028BF29BF028028BF57FC001528BF02800015288028BF500129BF;
defparam sp_inst_33.INIT_RAM_17 = 256'h57FB0280500129BF028028BF29BF028028BF57FC001528BF02800015288028BF;
defparam sp_inst_33.INIT_RAM_18 = 256'h001028BF028028BF001C028028BF500029BF29BF028028BF500129BF028028BF;
defparam sp_inst_33.INIT_RAM_19 = 256'h028028BF67FD02802800001028BF028028BF29BF028028BF29BF001002BF2800;
defparam sp_inst_33.INIT_RAM_1A = 256'h2800001028BF028028BF001C028028BF500029BF53FD67FF02802800001028BF;
defparam sp_inst_33.INIT_RAM_1B = 256'h28BF028028BF67FD02802800001028BF028028BF29BF028028BF29BF001002BF;
defparam sp_inst_33.INIT_RAM_1C = 256'h00152A3F57FA02805C000280283F5000034057FA028053FD67FF028028000010;
defparam sp_inst_33.INIT_RAM_1D = 256'h02BF4C000281288028800015001547FC2800001028BF28BF29BF028028BF57FA;
defparam sp_inst_33.INIT_RAM_1E = 256'h2880034029002A3F28BF43FF034000672A0028BF0340293F001529BF02802980;
defparam sp_inst_33.INIT_RAM_1F = 256'h0280298002BF4C0002802880034029800396154A157F0280298002BF4C000280;
defparam sp_inst_33.INIT_RAM_20 = 256'h00150014001728BF02802881157F440028BF29BF28BF6000028028BF29BF29BF;
defparam sp_inst_33.INIT_RAM_21 = 256'h02BF28BF500029810015157F0015001728BF02802881157F500029810014157F;
defparam sp_inst_33.INIT_RAM_22 = 256'h2881157F500029810014157F00150014001728BF02802881157F440028BF29BF;
defparam sp_inst_33.INIT_RAM_23 = 256'h29BF29BF0280298002BF4C0002802880034029810015157F0015001728BF0280;
defparam sp_inst_33.INIT_RAM_24 = 256'h0014157F00150014001728BF02802881157F440028BF29BF28BF6000028028BF;
defparam sp_inst_33.INIT_RAM_25 = 256'h28BF29BF02BF28BF500029810015157F0015001728BF02802881157F50002981;
defparam sp_inst_33.INIT_RAM_26 = 256'h28BF02802881157F500029810014157F00150014001728BF02802881157F4400;
defparam sp_inst_33.INIT_RAM_27 = 256'h2880157F29BF29BF0280298002BF4C0002802880034029810015157F00150017;
defparam sp_inst_33.INIT_RAM_28 = 256'h29BF0280298002BF4C0002802880001528BF29BF500029BF02804000001428BF;
defparam sp_inst_33.INIT_RAM_29 = 256'h03402900006703800380157F00672A000380157F2980001528BF157F2880157F;
defparam sp_inst_33.INIT_RAM_2A = 256'h1CC700152A3F2980028002951CC7293F001502802980298002BF4C0002802880;
defparam sp_inst_33.INIT_RAM_2B = 256'h28BF288028BF293F001529BF0280298002BF4C00028028802880034054000295;
defparam sp_inst_33.INIT_RAM_2C = 256'h298028BF6000288028BF288028BF298028BF0280288028BF29002A3F00102880;
defparam sp_inst_33.INIT_RAM_2D = 256'h288028BF298028BF288028BF6400288028BF288028BF298028BF0280288028BF;
defparam sp_inst_33.INIT_RAM_2E = 256'h298002BF4C00028028800340298028BF6000288028BF288028BF298028BF0280;
defparam sp_inst_33.INIT_RAM_2F = 256'h028057FB0280028057FC0280028057FC0280028057FC0280028057F502802980;
defparam sp_inst_33.INIT_RAM_30 = 256'h0280028057FB0280028057FB0280028057FB0280028057FB0280028057FB0280;
defparam sp_inst_33.INIT_RAM_31 = 256'h28BF0340034003400340500029BF03BF140057FB0280028057FB0280028057FB;
defparam sp_inst_33.INIT_RAM_32 = 256'h028057FC0280028057FC0280028057FC0280028057FC0280028047FF29BF02BF;
defparam sp_inst_33.INIT_RAM_33 = 256'h0280028057FB0280028057FC0280028057FC0280028057FC0280028057FC0280;
defparam sp_inst_33.INIT_RAM_34 = 256'h28BF0340034003400340500029BF03BF140057FB0280028057FB0280028057FB;
defparam sp_inst_33.INIT_RAM_35 = 256'h001557FB0280001557FB0280001557FB0280001557FB0280001547FF29BF02BF;
defparam sp_inst_33.INIT_RAM_36 = 256'h0280001557FB0280001557FB0280001557FB0280001557FB0280001557FB0280;
defparam sp_inst_33.INIT_RAM_37 = 256'h28BF0340034003400340500029BF03BF140057FB0280001557FB0280001557FB;
defparam sp_inst_33.INIT_RAM_38 = 256'h157F028057F502BA1C00028002811C0002802980298002BF53FE47FF29BF02BF;
defparam sp_inst_33.INIT_RAM_39 = 256'h02B81C00028002801C0002802980298002BF4C00028028802880034057F30380;
defparam sp_inst_33.INIT_RAM_3A = 256'h02801C0002802980298002BF4C00028028802880034057F30380157F028057F5;
defparam sp_inst_33.INIT_RAM_3B = 256'h2980298002BF4C00028028802880034057F20380157F028057F502B71C000280;
defparam sp_inst_33.INIT_RAM_3C = 256'h4C00028028802880034057F20380157F028057F402B61C00028002BF1C000280;
defparam sp_inst_33.INIT_RAM_3D = 256'h2880034057F20380157F028057F402B51C00028002BE1C0002802980298002BF;
defparam sp_inst_33.INIT_RAM_3E = 256'h0380157F028057F402B41C00028002BD1C0002802980298002BF4C0002802880;
defparam sp_inst_33.INIT_RAM_3F = 256'h57F302B31C00028002BC1C0002802980298002BF4C00028028802880034057F1;

SP sp_inst_34 (
    .DO({sp_inst_34_dout_w[15:0],sp_inst_34_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_2}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_34.READ_MODE = 1'b0;
defparam sp_inst_34.WRITE_MODE = 2'b01;
defparam sp_inst_34.BIT_WIDTH = 16;
defparam sp_inst_34.BLK_SEL = 3'b001;
defparam sp_inst_34.RESET_MODE = "SYNC";
defparam sp_inst_34.INIT_RAM_00 = 256'h028002BB1C0002802980298002BF4C00028028802880034057F10380157F0281;
defparam sp_inst_34.INIT_RAM_01 = 256'h02802980298002BF4C00028028802880034057F10380157F028257F302B11C00;
defparam sp_inst_34.INIT_RAM_02 = 256'h02BF4C00028028802880034057F00380157F028457F302B01C00028002BB1C00;
defparam sp_inst_34.INIT_RAM_03 = 256'h28802880034057F00380157F028857F202AF1C00028102BA1C00028029802980;
defparam sp_inst_34.INIT_RAM_04 = 256'h57F00380157F029057F202AE1C00028102B91C0002802980298002BF4C000280;
defparam sp_inst_34.INIT_RAM_05 = 256'h03A057F202AD1C00028102B81C0002802980298002BF4C000280288028800340;
defparam sp_inst_34.INIT_RAM_06 = 256'h1C00028102B71C0002802980298002BF4C00028028802880034057F00380157F;
defparam sp_inst_34.INIT_RAM_07 = 256'h1C0002802980298002BF4C00028028802880034057EF0380157F140057F202AB;
defparam sp_inst_34.INIT_RAM_08 = 256'h298002BF4C00028028802880034057EF0380157F140057F102AA1C00028102B7;
defparam sp_inst_34.INIT_RAM_09 = 256'h028028802880034057EF0380157F140057F102A91C00028102B61C0002802980;
defparam sp_inst_34.INIT_RAM_0A = 256'h034057EE0380157F140057F102A81C00028102B51C0002802980298002BF4C00;
defparam sp_inst_34.INIT_RAM_0B = 256'h157F140057F002A71C00028102B41C0002802980298002BF4C00028028802880;
defparam sp_inst_34.INIT_RAM_0C = 256'h02A51C00028102B31C0002802980298002BF4C00028028802880034057EE0380;
defparam sp_inst_34.INIT_RAM_0D = 256'h02B31C0002802980298002BF4C00028028802880034057EE0380157F140057F0;
defparam sp_inst_34.INIT_RAM_0E = 256'h2980298002BF4C00028028802880034057ED0380157F140057F002A41C000281;
defparam sp_inst_34.INIT_RAM_0F = 256'h4C00028028802880034057ED0380157F140057F002A31C00028102B21C000280;
defparam sp_inst_34.INIT_RAM_10 = 256'h2880034057ED0380157F140057EF02A21C00028202B11C0002802980298002BF;
defparam sp_inst_34.INIT_RAM_11 = 256'h0380157F140057EF02A11C00028202B01C0002802980298002BF4C0002802880;
defparam sp_inst_34.INIT_RAM_12 = 256'h57EF02A01C00028202AF1C0002802980298002BF4C00028028802880034057ED;
defparam sp_inst_34.INIT_RAM_13 = 256'h028202AE1C0002802980298002BF4C00028028802880034057EC0380157F1400;
defparam sp_inst_34.INIT_RAM_14 = 256'h02802980298002BF4C00028028802880034057EC0380157F140157EE029E1C00;
defparam sp_inst_34.INIT_RAM_15 = 256'h02BF4C00028028802880034057EC0380157F140257EE029D1C00028202AE1C00;
defparam sp_inst_34.INIT_RAM_16 = 256'h28802880034057EB0380157F140457EE029C1C00028202AD1C00028029802980;
defparam sp_inst_34.INIT_RAM_17 = 256'h57EB0380157F140857ED029B1C00028202AC1C0002802980298002BF4C000280;
defparam sp_inst_34.INIT_RAM_18 = 256'h141057ED029A1C00028202AB1C0002802980298002BF4C000280288028800340;
defparam sp_inst_34.INIT_RAM_19 = 256'h1C00028202AA1C0002802980298002BF4C00028028802880034057EB0380157F;
defparam sp_inst_34.INIT_RAM_1A = 256'h1C0002802980298002BF4C00028028802880034057EA0380157F142057ED0298;
defparam sp_inst_34.INIT_RAM_1B = 256'h298002BF4C00028028802880034057EA0380157F144057ED02971C00028202AA;
defparam sp_inst_34.INIT_RAM_1C = 256'h028028802880034057EA0380157F148057EC02961C00028202A91C0002802980;
defparam sp_inst_34.INIT_RAM_1D = 256'h034057EA0380157F150057EC02951C00028302A81C0002802980298002BF4C00;
defparam sp_inst_34.INIT_RAM_1E = 256'h1C00028302A71C00298014020380157F02802980298002BF4C00028028802880;
defparam sp_inst_34.INIT_RAM_1F = 256'h29BF034029BF001428BF28BF29BF28800380157F29BF28800380157F57EC0293;
defparam sp_inst_34.INIT_RAM_20 = 256'h29BF028028BF4C0028800010004028BF02961C0040000340001728BF28BF5000;
defparam sp_inst_34.INIT_RAM_21 = 256'h298014000380157F02802980298002BF4C0002802880288003406FFF028028BF;
defparam sp_inst_34.INIT_RAM_22 = 256'h0380157F02802980298002BF4C00028028802880034057EF29BF28800380157F;
defparam sp_inst_34.INIT_RAM_23 = 256'h157F298014000380157F293F0340006728800380157F297F037F006F00442880;
defparam sp_inst_34.INIT_RAM_24 = 256'h0280298002BF4C00028028802880034057EA028F1C0000152A7F298002800380;
defparam sp_inst_34.INIT_RAM_25 = 256'h02802980298002BF4C00028028800340293F2A000380157F298014000380157F;
defparam sp_inst_34.INIT_RAM_26 = 256'h028028BF2980001414010380157F28800380157F29BF0340004428800380157F;
defparam sp_inst_34.INIT_RAM_27 = 256'h1C00500029800380157F57E9028C1C004C002880001002911C00004028BF6800;
defparam sp_inst_34.INIT_RAM_28 = 256'h288028800340034050002980001403BF15FF0380157F28800380157F57E9028D;
defparam sp_inst_34.INIT_RAM_29 = 256'h001557EF0284400003402A3F293F2A000380157F02802980298002BF4C000280;
defparam sp_inst_34.INIT_RAM_2A = 256'h028B1C0000152A3F293F2A00157F400003402A3F57E9028B1C0057EF02844000;
defparam sp_inst_34.INIT_RAM_2B = 256'h0380157F57EF00152A3F293F2A00157F400003402A3F290002800380157F57E9;
defparam sp_inst_34.INIT_RAM_2C = 256'h57E602802980298002BF4C000280288028800340290002BF0380157F29000280;
defparam sp_inst_34.INIT_RAM_2D = 256'h1C001C001C001C001C001C001C004C00028028802880034057E657E802891C00;
defparam sp_inst_34.INIT_RAM_2E = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_34.INIT_RAM_2F = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_34.INIT_RAM_30 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_34.INIT_RAM_31 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_34.INIT_RAM_32 = 256'h203A696C3C201C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_34.INIT_RAM_33 = 256'h2D2D00002E2E2E2E2E2E2E2E495F4F532E2E2E2E2E2E00000A0D20203A636620;
defparam sp_inst_34.INIT_RAM_34 = 256'h2E2E2E2E2E2E2E2E414641422E2E2E2E2E2E000078253A6C6E617965746E6375;
defparam sp_inst_34.INIT_RAM_35 = 256'h20726C63656D20737265697200000A2E2E2E2E2E2E2E44412E2E2E2E2E2E0000;
defparam sp_inst_34.INIT_RAM_36 = 256'h2E2E7572746E726163206D69657200000A78303A6572747200000A2E70756574;
defparam sp_inst_34.INIT_RAM_37 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C000000;
defparam sp_inst_34.INIT_RAM_38 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_34.INIT_RAM_39 = 256'h1C001C001C001C001C001C001C001C001C001C001C001C001C001C001C001C00;
defparam sp_inst_34.INIT_RAM_3A = 256'h697069740072646E5F715F31697069740072646E5F715F30697069741C001C00;
defparam sp_inst_34.INIT_RAM_3B = 256'h0072646E5F715F34697069740072646E5F715F33697069740072646E5F715F32;
defparam sp_inst_34.INIT_RAM_3C = 256'h5F715F37697069740072646E5F715F36697069740072646E5F715F3569706974;
defparam sp_inst_34.INIT_RAM_3D = 256'h697069740072646E5F715F31697069740072646E5F715F30697069740072646E;
defparam sp_inst_34.INIT_RAM_3E = 256'h0072646E5F715F34697069740072646E5F715F33697069740072646E5F715F32;
defparam sp_inst_34.INIT_RAM_3F = 256'h5F715F37697069740072646E5F715F36697069740072646E5F715F3569706974;

SP sp_inst_35 (
    .DO({sp_inst_35_dout_w[15:0],sp_inst_35_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_3}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_35.READ_MODE = 1'b0;
defparam sp_inst_35.WRITE_MODE = 2'b01;
defparam sp_inst_35.BIT_WIDTH = 16;
defparam sp_inst_35.BLK_SEL = 3'b001;
defparam sp_inst_35.RESET_MODE = "SYNC";
defparam sp_inst_35.INIT_RAM_00 = 256'h697069740072646E5F715F31697069740072646E5F715F30697069740072646E;
defparam sp_inst_35.INIT_RAM_01 = 256'h0072646E5F715F34697069740072646E5F715F33697069740072646E5F715F32;
defparam sp_inst_35.INIT_RAM_02 = 256'h5F715F37697069740072646E5F715F36697069740072646E5F715F3569706974;
defparam sp_inst_35.INIT_RAM_03 = 256'h697069740072646E5F715F31697069740072646E5F715F30697069740072646E;
defparam sp_inst_35.INIT_RAM_04 = 256'h0072646E5F715F34697069740072646E5F715F33697069740072646E5F715F32;
defparam sp_inst_35.INIT_RAM_05 = 256'h5F715F37697069740072646E5F715F36697069740072646E5F715F3569706974;
defparam sp_inst_35.INIT_RAM_06 = 256'h000000000000000000000000000000000000000000000072646E5F740072646E;
defparam sp_inst_35.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_35.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_36 (
    .DO({sp_inst_36_dout_w[15:0],sp_inst_36_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_4}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_36.READ_MODE = 1'b0;
defparam sp_inst_36.WRITE_MODE = 2'b01;
defparam sp_inst_36.BIT_WIDTH = 16;
defparam sp_inst_36.BLK_SEL = 3'b001;
defparam sp_inst_36.RESET_MODE = "SYNC";
defparam sp_inst_36.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_36.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_37 (
    .DO({sp_inst_37_dout_w[15:0],sp_inst_37_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_5}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_37.READ_MODE = 1'b0;
defparam sp_inst_37.WRITE_MODE = 2'b01;
defparam sp_inst_37.BIT_WIDTH = 16;
defparam sp_inst_37.BLK_SEL = 3'b001;
defparam sp_inst_37.RESET_MODE = "SYNC";
defparam sp_inst_37.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_37.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_38 (
    .DO({sp_inst_38_dout_w[15:0],sp_inst_38_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_6}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_38.READ_MODE = 1'b0;
defparam sp_inst_38.WRITE_MODE = 2'b01;
defparam sp_inst_38.BIT_WIDTH = 16;
defparam sp_inst_38.BLK_SEL = 3'b001;
defparam sp_inst_38.RESET_MODE = "SYNC";
defparam sp_inst_38.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_38.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_39 (
    .DO({sp_inst_39_dout_w[15:0],sp_inst_39_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_7}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_39.READ_MODE = 1'b0;
defparam sp_inst_39.WRITE_MODE = 2'b01;
defparam sp_inst_39.BIT_WIDTH = 16;
defparam sp_inst_39.BLK_SEL = 3'b001;
defparam sp_inst_39.RESET_MODE = "SYNC";
defparam sp_inst_39.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_39.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_40 (
    .DO({sp_inst_40_dout_w[15:0],sp_inst_40_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_8}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_40.READ_MODE = 1'b0;
defparam sp_inst_40.WRITE_MODE = 2'b01;
defparam sp_inst_40.BIT_WIDTH = 16;
defparam sp_inst_40.BLK_SEL = 3'b001;
defparam sp_inst_40.RESET_MODE = "SYNC";
defparam sp_inst_40.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_40.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_41 (
    .DO({sp_inst_41_dout_w[15:0],sp_inst_41_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_9}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_41.READ_MODE = 1'b0;
defparam sp_inst_41.WRITE_MODE = 2'b01;
defparam sp_inst_41.BIT_WIDTH = 16;
defparam sp_inst_41.BLK_SEL = 3'b001;
defparam sp_inst_41.RESET_MODE = "SYNC";
defparam sp_inst_41.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_41.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_42 (
    .DO({sp_inst_42_dout_w[15:0],sp_inst_42_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_10}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_42.READ_MODE = 1'b0;
defparam sp_inst_42.WRITE_MODE = 2'b01;
defparam sp_inst_42.BIT_WIDTH = 16;
defparam sp_inst_42.BLK_SEL = 3'b001;
defparam sp_inst_42.RESET_MODE = "SYNC";
defparam sp_inst_42.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_42.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_43 (
    .DO({sp_inst_43_dout_w[15:0],sp_inst_43_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_11}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_43.READ_MODE = 1'b0;
defparam sp_inst_43.WRITE_MODE = 2'b01;
defparam sp_inst_43.BIT_WIDTH = 16;
defparam sp_inst_43.BLK_SEL = 3'b001;
defparam sp_inst_43.RESET_MODE = "SYNC";
defparam sp_inst_43.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_43.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_44 (
    .DO({sp_inst_44_dout_w[15:0],sp_inst_44_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_12}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_44.READ_MODE = 1'b0;
defparam sp_inst_44.WRITE_MODE = 2'b01;
defparam sp_inst_44.BIT_WIDTH = 16;
defparam sp_inst_44.BLK_SEL = 3'b001;
defparam sp_inst_44.RESET_MODE = "SYNC";
defparam sp_inst_44.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_44.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_45 (
    .DO({sp_inst_45_dout_w[15:0],sp_inst_45_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_13}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_45.READ_MODE = 1'b0;
defparam sp_inst_45.WRITE_MODE = 2'b01;
defparam sp_inst_45.BIT_WIDTH = 16;
defparam sp_inst_45.BLK_SEL = 3'b001;
defparam sp_inst_45.RESET_MODE = "SYNC";
defparam sp_inst_45.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_45.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_46 (
    .DO({sp_inst_46_dout_w[15:0],sp_inst_46_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_14}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_46.READ_MODE = 1'b0;
defparam sp_inst_46.WRITE_MODE = 2'b01;
defparam sp_inst_46.BIT_WIDTH = 16;
defparam sp_inst_46.BLK_SEL = 3'b001;
defparam sp_inst_46.RESET_MODE = "SYNC";
defparam sp_inst_46.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_46.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_47 (
    .DO({sp_inst_47_dout_w[15:0],sp_inst_47_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_15}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_47.READ_MODE = 1'b0;
defparam sp_inst_47.WRITE_MODE = 2'b01;
defparam sp_inst_47.BIT_WIDTH = 16;
defparam sp_inst_47.BLK_SEL = 3'b001;
defparam sp_inst_47.RESET_MODE = "SYNC";
defparam sp_inst_47.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_47.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_48 (
    .DO({sp_inst_48_dout_w[15:0],sp_inst_48_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_16}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_48.READ_MODE = 1'b0;
defparam sp_inst_48.WRITE_MODE = 2'b01;
defparam sp_inst_48.BIT_WIDTH = 16;
defparam sp_inst_48.BLK_SEL = 3'b001;
defparam sp_inst_48.RESET_MODE = "SYNC";
defparam sp_inst_48.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_48.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_49 (
    .DO({sp_inst_49_dout_w[15:0],sp_inst_49_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_17}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_49.READ_MODE = 1'b0;
defparam sp_inst_49.WRITE_MODE = 2'b01;
defparam sp_inst_49.BIT_WIDTH = 16;
defparam sp_inst_49.BLK_SEL = 3'b001;
defparam sp_inst_49.RESET_MODE = "SYNC";
defparam sp_inst_49.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_49.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_50 (
    .DO({sp_inst_50_dout_w[15:0],sp_inst_50_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_18}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_50.READ_MODE = 1'b0;
defparam sp_inst_50.WRITE_MODE = 2'b01;
defparam sp_inst_50.BIT_WIDTH = 16;
defparam sp_inst_50.BLK_SEL = 3'b001;
defparam sp_inst_50.RESET_MODE = "SYNC";
defparam sp_inst_50.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_50.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_51 (
    .DO({sp_inst_51_dout_w[15:0],sp_inst_51_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_19}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_51.READ_MODE = 1'b0;
defparam sp_inst_51.WRITE_MODE = 2'b01;
defparam sp_inst_51.BIT_WIDTH = 16;
defparam sp_inst_51.BLK_SEL = 3'b001;
defparam sp_inst_51.RESET_MODE = "SYNC";
defparam sp_inst_51.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_51.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_52 (
    .DO({sp_inst_52_dout_w[15:0],sp_inst_52_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_20}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_52.READ_MODE = 1'b0;
defparam sp_inst_52.WRITE_MODE = 2'b01;
defparam sp_inst_52.BIT_WIDTH = 16;
defparam sp_inst_52.BLK_SEL = 3'b001;
defparam sp_inst_52.RESET_MODE = "SYNC";
defparam sp_inst_52.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_52.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_53 (
    .DO({sp_inst_53_dout_w[15:0],sp_inst_53_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_21}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_53.READ_MODE = 1'b0;
defparam sp_inst_53.WRITE_MODE = 2'b01;
defparam sp_inst_53.BIT_WIDTH = 16;
defparam sp_inst_53.BLK_SEL = 3'b001;
defparam sp_inst_53.RESET_MODE = "SYNC";
defparam sp_inst_53.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_53.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_54 (
    .DO({sp_inst_54_dout_w[15:0],sp_inst_54_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_22}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_54.READ_MODE = 1'b0;
defparam sp_inst_54.WRITE_MODE = 2'b01;
defparam sp_inst_54.BIT_WIDTH = 16;
defparam sp_inst_54.BLK_SEL = 3'b001;
defparam sp_inst_54.RESET_MODE = "SYNC";
defparam sp_inst_54.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_54.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_55 (
    .DO({sp_inst_55_dout_w[15:0],sp_inst_55_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_23}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_55.READ_MODE = 1'b0;
defparam sp_inst_55.WRITE_MODE = 2'b01;
defparam sp_inst_55.BIT_WIDTH = 16;
defparam sp_inst_55.BLK_SEL = 3'b001;
defparam sp_inst_55.RESET_MODE = "SYNC";
defparam sp_inst_55.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_55.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_56 (
    .DO({sp_inst_56_dout_w[15:0],sp_inst_56_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_24}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_56.READ_MODE = 1'b0;
defparam sp_inst_56.WRITE_MODE = 2'b01;
defparam sp_inst_56.BIT_WIDTH = 16;
defparam sp_inst_56.BLK_SEL = 3'b001;
defparam sp_inst_56.RESET_MODE = "SYNC";
defparam sp_inst_56.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_56.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_57 (
    .DO({sp_inst_57_dout_w[15:0],sp_inst_57_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_25}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_57.READ_MODE = 1'b0;
defparam sp_inst_57.WRITE_MODE = 2'b01;
defparam sp_inst_57.BIT_WIDTH = 16;
defparam sp_inst_57.BLK_SEL = 3'b001;
defparam sp_inst_57.RESET_MODE = "SYNC";
defparam sp_inst_57.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_57.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_58 (
    .DO({sp_inst_58_dout_w[15:0],sp_inst_58_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_26}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_58.READ_MODE = 1'b0;
defparam sp_inst_58.WRITE_MODE = 2'b01;
defparam sp_inst_58.BIT_WIDTH = 16;
defparam sp_inst_58.BLK_SEL = 3'b001;
defparam sp_inst_58.RESET_MODE = "SYNC";
defparam sp_inst_58.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_58.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_59 (
    .DO({sp_inst_59_dout_w[15:0],sp_inst_59_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_27}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_59.READ_MODE = 1'b0;
defparam sp_inst_59.WRITE_MODE = 2'b01;
defparam sp_inst_59.BIT_WIDTH = 16;
defparam sp_inst_59.BLK_SEL = 3'b001;
defparam sp_inst_59.RESET_MODE = "SYNC";
defparam sp_inst_59.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_59.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_60 (
    .DO({sp_inst_60_dout_w[15:0],sp_inst_60_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_28}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_60.READ_MODE = 1'b0;
defparam sp_inst_60.WRITE_MODE = 2'b01;
defparam sp_inst_60.BIT_WIDTH = 16;
defparam sp_inst_60.BLK_SEL = 3'b001;
defparam sp_inst_60.RESET_MODE = "SYNC";
defparam sp_inst_60.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_60.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_61 (
    .DO({sp_inst_61_dout_w[15:0],sp_inst_61_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_29}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_61.READ_MODE = 1'b0;
defparam sp_inst_61.WRITE_MODE = 2'b01;
defparam sp_inst_61.BIT_WIDTH = 16;
defparam sp_inst_61.BLK_SEL = 3'b001;
defparam sp_inst_61.RESET_MODE = "SYNC";
defparam sp_inst_61.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_61.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_62 (
    .DO({sp_inst_62_dout_w[15:0],sp_inst_62_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_30}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_62.READ_MODE = 1'b0;
defparam sp_inst_62.WRITE_MODE = 2'b01;
defparam sp_inst_62.BIT_WIDTH = 16;
defparam sp_inst_62.BLK_SEL = 3'b001;
defparam sp_inst_62.RESET_MODE = "SYNC";
defparam sp_inst_62.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_62.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_63 (
    .DO({sp_inst_63_dout_w[15:0],sp_inst_63_dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_31}),
    .AD({ad[9:0],gw_gnd,gw_gnd,byte_en[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_63.READ_MODE = 1'b0;
defparam sp_inst_63.WRITE_MODE = 2'b01;
defparam sp_inst_63.BIT_WIDTH = 16;
defparam sp_inst_63.BLK_SEL = 3'b001;
defparam sp_inst_63.RESET_MODE = "SYNC";
defparam sp_inst_63.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_63.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
DFFRE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
DFFRE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
DFFRE dff_inst_3 (
  .Q(dff_q_3),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
DFFRE dff_inst_4 (
  .Q(dff_q_4),
  .D(ad[10]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(sp_inst_0_dout[0]),
  .I1(sp_inst_1_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(sp_inst_2_dout[0]),
  .I1(sp_inst_3_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(sp_inst_4_dout[0]),
  .I1(sp_inst_5_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(sp_inst_6_dout[0]),
  .I1(sp_inst_7_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(sp_inst_8_dout[0]),
  .I1(sp_inst_9_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(sp_inst_10_dout[0]),
  .I1(sp_inst_11_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(sp_inst_12_dout[0]),
  .I1(sp_inst_13_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(sp_inst_14_dout[0]),
  .I1(sp_inst_15_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(sp_inst_16_dout[0]),
  .I1(sp_inst_17_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(sp_inst_18_dout[0]),
  .I1(sp_inst_19_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(sp_inst_20_dout[0]),
  .I1(sp_inst_21_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(sp_inst_22_dout[0]),
  .I1(sp_inst_23_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(sp_inst_24_dout[0]),
  .I1(sp_inst_25_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(sp_inst_26_dout[0]),
  .I1(sp_inst_27_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(sp_inst_28_dout[0]),
  .I1(sp_inst_29_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(sp_inst_30_dout[0]),
  .I1(sp_inst_31_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_3)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_3)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_3)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(dff_q_3)
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(dff_q_3)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_3)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_3)
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(dff_q_3)
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(dff_q_2)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(dff_q_2)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(mux_o_20),
  .I1(mux_o_21),
  .S0(dff_q_2)
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(mux_o_22),
  .I1(mux_o_23),
  .S0(dff_q_2)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(mux_o_24),
  .I1(mux_o_25),
  .S0(dff_q_1)
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(mux_o_26),
  .I1(mux_o_27),
  .S0(dff_q_1)
);
MUX2 mux_inst_30 (
  .O(dout[0]),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(dff_q_0)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(sp_inst_0_dout[1]),
  .I1(sp_inst_1_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(sp_inst_2_dout[1]),
  .I1(sp_inst_3_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(sp_inst_4_dout[1]),
  .I1(sp_inst_5_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(sp_inst_6_dout[1]),
  .I1(sp_inst_7_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(sp_inst_8_dout[1]),
  .I1(sp_inst_9_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(sp_inst_10_dout[1]),
  .I1(sp_inst_11_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(sp_inst_12_dout[1]),
  .I1(sp_inst_13_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(sp_inst_14_dout[1]),
  .I1(sp_inst_15_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(sp_inst_16_dout[1]),
  .I1(sp_inst_17_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(sp_inst_18_dout[1]),
  .I1(sp_inst_19_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(sp_inst_20_dout[1]),
  .I1(sp_inst_21_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(sp_inst_22_dout[1]),
  .I1(sp_inst_23_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(sp_inst_24_dout[1]),
  .I1(sp_inst_25_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(sp_inst_26_dout[1]),
  .I1(sp_inst_27_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(sp_inst_28_dout[1]),
  .I1(sp_inst_29_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(sp_inst_30_dout[1]),
  .I1(sp_inst_31_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(mux_o_31),
  .I1(mux_o_32),
  .S0(dff_q_3)
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(mux_o_33),
  .I1(mux_o_34),
  .S0(dff_q_3)
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(mux_o_35),
  .I1(mux_o_36),
  .S0(dff_q_3)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(mux_o_37),
  .I1(mux_o_38),
  .S0(dff_q_3)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(mux_o_39),
  .I1(mux_o_40),
  .S0(dff_q_3)
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(mux_o_41),
  .I1(mux_o_42),
  .S0(dff_q_3)
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_43),
  .I1(mux_o_44),
  .S0(dff_q_3)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(dff_q_3)
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(mux_o_47),
  .I1(mux_o_48),
  .S0(dff_q_2)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(dff_q_2)
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(mux_o_51),
  .I1(mux_o_52),
  .S0(dff_q_2)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(mux_o_53),
  .I1(mux_o_54),
  .S0(dff_q_2)
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(mux_o_55),
  .I1(mux_o_56),
  .S0(dff_q_1)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(mux_o_57),
  .I1(mux_o_58),
  .S0(dff_q_1)
);
MUX2 mux_inst_61 (
  .O(dout[1]),
  .I0(mux_o_59),
  .I1(mux_o_60),
  .S0(dff_q_0)
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(sp_inst_0_dout[2]),
  .I1(sp_inst_1_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(sp_inst_2_dout[2]),
  .I1(sp_inst_3_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(sp_inst_4_dout[2]),
  .I1(sp_inst_5_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(sp_inst_6_dout[2]),
  .I1(sp_inst_7_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(sp_inst_8_dout[2]),
  .I1(sp_inst_9_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(sp_inst_10_dout[2]),
  .I1(sp_inst_11_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(sp_inst_12_dout[2]),
  .I1(sp_inst_13_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(sp_inst_14_dout[2]),
  .I1(sp_inst_15_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(sp_inst_16_dout[2]),
  .I1(sp_inst_17_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(sp_inst_18_dout[2]),
  .I1(sp_inst_19_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(sp_inst_20_dout[2]),
  .I1(sp_inst_21_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(sp_inst_22_dout[2]),
  .I1(sp_inst_23_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(sp_inst_24_dout[2]),
  .I1(sp_inst_25_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(sp_inst_26_dout[2]),
  .I1(sp_inst_27_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(sp_inst_28_dout[2]),
  .I1(sp_inst_29_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(sp_inst_30_dout[2]),
  .I1(sp_inst_31_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(dff_q_3)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(mux_o_64),
  .I1(mux_o_65),
  .S0(dff_q_3)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(dff_q_3)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(mux_o_68),
  .I1(mux_o_69),
  .S0(dff_q_3)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(dff_q_3)
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(dff_q_3)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(mux_o_74),
  .I1(mux_o_75),
  .S0(dff_q_3)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(mux_o_76),
  .I1(mux_o_77),
  .S0(dff_q_3)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(mux_o_78),
  .I1(mux_o_79),
  .S0(dff_q_2)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(mux_o_80),
  .I1(mux_o_81),
  .S0(dff_q_2)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_82),
  .I1(mux_o_83),
  .S0(dff_q_2)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(mux_o_84),
  .I1(mux_o_85),
  .S0(dff_q_2)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(mux_o_86),
  .I1(mux_o_87),
  .S0(dff_q_1)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(mux_o_88),
  .I1(mux_o_89),
  .S0(dff_q_1)
);
MUX2 mux_inst_92 (
  .O(dout[2]),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(dff_q_0)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(sp_inst_0_dout[3]),
  .I1(sp_inst_1_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(sp_inst_2_dout[3]),
  .I1(sp_inst_3_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(sp_inst_4_dout[3]),
  .I1(sp_inst_5_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(sp_inst_6_dout[3]),
  .I1(sp_inst_7_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(sp_inst_8_dout[3]),
  .I1(sp_inst_9_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(sp_inst_10_dout[3]),
  .I1(sp_inst_11_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(sp_inst_12_dout[3]),
  .I1(sp_inst_13_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(sp_inst_14_dout[3]),
  .I1(sp_inst_15_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(sp_inst_16_dout[3]),
  .I1(sp_inst_17_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(sp_inst_18_dout[3]),
  .I1(sp_inst_19_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(sp_inst_20_dout[3]),
  .I1(sp_inst_21_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_104 (
  .O(mux_o_104),
  .I0(sp_inst_22_dout[3]),
  .I1(sp_inst_23_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(sp_inst_24_dout[3]),
  .I1(sp_inst_25_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(sp_inst_26_dout[3]),
  .I1(sp_inst_27_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(sp_inst_28_dout[3]),
  .I1(sp_inst_29_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(sp_inst_30_dout[3]),
  .I1(sp_inst_31_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(mux_o_93),
  .I1(mux_o_94),
  .S0(dff_q_3)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(mux_o_95),
  .I1(mux_o_96),
  .S0(dff_q_3)
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(mux_o_97),
  .I1(mux_o_98),
  .S0(dff_q_3)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(mux_o_99),
  .I1(mux_o_100),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_101),
  .I1(mux_o_102),
  .S0(dff_q_3)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_103),
  .I1(mux_o_104),
  .S0(dff_q_3)
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(dff_q_3)
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(dff_q_3)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(dff_q_2)
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_111),
  .I1(mux_o_112),
  .S0(dff_q_2)
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(mux_o_113),
  .I1(mux_o_114),
  .S0(dff_q_2)
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(mux_o_115),
  .I1(mux_o_116),
  .S0(dff_q_2)
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(mux_o_117),
  .I1(mux_o_118),
  .S0(dff_q_1)
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(mux_o_119),
  .I1(mux_o_120),
  .S0(dff_q_1)
);
MUX2 mux_inst_123 (
  .O(dout[3]),
  .I0(mux_o_121),
  .I1(mux_o_122),
  .S0(dff_q_0)
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(sp_inst_0_dout[4]),
  .I1(sp_inst_1_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_125 (
  .O(mux_o_125),
  .I0(sp_inst_2_dout[4]),
  .I1(sp_inst_3_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(sp_inst_4_dout[4]),
  .I1(sp_inst_5_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(sp_inst_6_dout[4]),
  .I1(sp_inst_7_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(sp_inst_8_dout[4]),
  .I1(sp_inst_9_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(sp_inst_10_dout[4]),
  .I1(sp_inst_11_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(sp_inst_12_dout[4]),
  .I1(sp_inst_13_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(sp_inst_14_dout[4]),
  .I1(sp_inst_15_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(sp_inst_16_dout[4]),
  .I1(sp_inst_17_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(sp_inst_18_dout[4]),
  .I1(sp_inst_19_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(sp_inst_20_dout[4]),
  .I1(sp_inst_21_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(sp_inst_22_dout[4]),
  .I1(sp_inst_23_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(sp_inst_24_dout[4]),
  .I1(sp_inst_25_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(sp_inst_26_dout[4]),
  .I1(sp_inst_27_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(sp_inst_28_dout[4]),
  .I1(sp_inst_29_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(sp_inst_30_dout[4]),
  .I1(sp_inst_31_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(mux_o_124),
  .I1(mux_o_125),
  .S0(dff_q_3)
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(dff_q_3)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(dff_q_3)
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(dff_q_3)
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(mux_o_132),
  .I1(mux_o_133),
  .S0(dff_q_3)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(mux_o_134),
  .I1(mux_o_135),
  .S0(dff_q_3)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(mux_o_136),
  .I1(mux_o_137),
  .S0(dff_q_3)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(mux_o_138),
  .I1(mux_o_139),
  .S0(dff_q_3)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(mux_o_140),
  .I1(mux_o_141),
  .S0(dff_q_2)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(mux_o_142),
  .I1(mux_o_143),
  .S0(dff_q_2)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(mux_o_144),
  .I1(mux_o_145),
  .S0(dff_q_2)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(mux_o_146),
  .I1(mux_o_147),
  .S0(dff_q_2)
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(mux_o_148),
  .I1(mux_o_149),
  .S0(dff_q_1)
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(mux_o_150),
  .I1(mux_o_151),
  .S0(dff_q_1)
);
MUX2 mux_inst_154 (
  .O(dout[4]),
  .I0(mux_o_152),
  .I1(mux_o_153),
  .S0(dff_q_0)
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(sp_inst_0_dout[5]),
  .I1(sp_inst_1_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(sp_inst_2_dout[5]),
  .I1(sp_inst_3_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(sp_inst_4_dout[5]),
  .I1(sp_inst_5_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(sp_inst_6_dout[5]),
  .I1(sp_inst_7_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(sp_inst_8_dout[5]),
  .I1(sp_inst_9_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(sp_inst_10_dout[5]),
  .I1(sp_inst_11_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(sp_inst_12_dout[5]),
  .I1(sp_inst_13_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(sp_inst_14_dout[5]),
  .I1(sp_inst_15_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(sp_inst_16_dout[5]),
  .I1(sp_inst_17_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(sp_inst_18_dout[5]),
  .I1(sp_inst_19_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(sp_inst_20_dout[5]),
  .I1(sp_inst_21_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(sp_inst_22_dout[5]),
  .I1(sp_inst_23_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(sp_inst_24_dout[5]),
  .I1(sp_inst_25_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(sp_inst_26_dout[5]),
  .I1(sp_inst_27_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(sp_inst_28_dout[5]),
  .I1(sp_inst_29_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(sp_inst_30_dout[5]),
  .I1(sp_inst_31_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(mux_o_155),
  .I1(mux_o_156),
  .S0(dff_q_3)
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(mux_o_157),
  .I1(mux_o_158),
  .S0(dff_q_3)
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(mux_o_159),
  .I1(mux_o_160),
  .S0(dff_q_3)
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(mux_o_161),
  .I1(mux_o_162),
  .S0(dff_q_3)
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(mux_o_163),
  .I1(mux_o_164),
  .S0(dff_q_3)
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(dff_q_3)
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(mux_o_167),
  .I1(mux_o_168),
  .S0(dff_q_3)
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(mux_o_169),
  .I1(mux_o_170),
  .S0(dff_q_3)
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(mux_o_171),
  .I1(mux_o_172),
  .S0(dff_q_2)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(mux_o_173),
  .I1(mux_o_174),
  .S0(dff_q_2)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(mux_o_175),
  .I1(mux_o_176),
  .S0(dff_q_2)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(mux_o_177),
  .I1(mux_o_178),
  .S0(dff_q_2)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(mux_o_179),
  .I1(mux_o_180),
  .S0(dff_q_1)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(mux_o_181),
  .I1(mux_o_182),
  .S0(dff_q_1)
);
MUX2 mux_inst_185 (
  .O(dout[5]),
  .I0(mux_o_183),
  .I1(mux_o_184),
  .S0(dff_q_0)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(sp_inst_0_dout[6]),
  .I1(sp_inst_1_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(sp_inst_2_dout[6]),
  .I1(sp_inst_3_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(sp_inst_4_dout[6]),
  .I1(sp_inst_5_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(sp_inst_6_dout[6]),
  .I1(sp_inst_7_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(sp_inst_8_dout[6]),
  .I1(sp_inst_9_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(sp_inst_10_dout[6]),
  .I1(sp_inst_11_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(sp_inst_12_dout[6]),
  .I1(sp_inst_13_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(sp_inst_14_dout[6]),
  .I1(sp_inst_15_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(sp_inst_16_dout[6]),
  .I1(sp_inst_17_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(sp_inst_18_dout[6]),
  .I1(sp_inst_19_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(sp_inst_20_dout[6]),
  .I1(sp_inst_21_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(sp_inst_22_dout[6]),
  .I1(sp_inst_23_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(sp_inst_24_dout[6]),
  .I1(sp_inst_25_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(sp_inst_26_dout[6]),
  .I1(sp_inst_27_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(sp_inst_28_dout[6]),
  .I1(sp_inst_29_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(sp_inst_30_dout[6]),
  .I1(sp_inst_31_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(dff_q_3)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_188),
  .I1(mux_o_189),
  .S0(dff_q_3)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(mux_o_190),
  .I1(mux_o_191),
  .S0(dff_q_3)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_192),
  .I1(mux_o_193),
  .S0(dff_q_3)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_194),
  .I1(mux_o_195),
  .S0(dff_q_3)
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(mux_o_196),
  .I1(mux_o_197),
  .S0(dff_q_3)
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(mux_o_198),
  .I1(mux_o_199),
  .S0(dff_q_3)
);
MUX2 mux_inst_209 (
  .O(mux_o_209),
  .I0(mux_o_200),
  .I1(mux_o_201),
  .S0(dff_q_3)
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(mux_o_202),
  .I1(mux_o_203),
  .S0(dff_q_2)
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(mux_o_204),
  .I1(mux_o_205),
  .S0(dff_q_2)
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(mux_o_206),
  .I1(mux_o_207),
  .S0(dff_q_2)
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(mux_o_208),
  .I1(mux_o_209),
  .S0(dff_q_2)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(mux_o_210),
  .I1(mux_o_211),
  .S0(dff_q_1)
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(mux_o_212),
  .I1(mux_o_213),
  .S0(dff_q_1)
);
MUX2 mux_inst_216 (
  .O(dout[6]),
  .I0(mux_o_214),
  .I1(mux_o_215),
  .S0(dff_q_0)
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(sp_inst_0_dout[7]),
  .I1(sp_inst_1_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(sp_inst_2_dout[7]),
  .I1(sp_inst_3_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(sp_inst_4_dout[7]),
  .I1(sp_inst_5_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(sp_inst_6_dout[7]),
  .I1(sp_inst_7_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(sp_inst_8_dout[7]),
  .I1(sp_inst_9_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(sp_inst_10_dout[7]),
  .I1(sp_inst_11_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(sp_inst_12_dout[7]),
  .I1(sp_inst_13_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(sp_inst_14_dout[7]),
  .I1(sp_inst_15_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(sp_inst_16_dout[7]),
  .I1(sp_inst_17_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(sp_inst_18_dout[7]),
  .I1(sp_inst_19_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(sp_inst_20_dout[7]),
  .I1(sp_inst_21_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(sp_inst_22_dout[7]),
  .I1(sp_inst_23_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(sp_inst_24_dout[7]),
  .I1(sp_inst_25_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(sp_inst_26_dout[7]),
  .I1(sp_inst_27_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(sp_inst_28_dout[7]),
  .I1(sp_inst_29_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(sp_inst_30_dout[7]),
  .I1(sp_inst_31_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_217),
  .I1(mux_o_218),
  .S0(dff_q_3)
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(mux_o_219),
  .I1(mux_o_220),
  .S0(dff_q_3)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_221),
  .I1(mux_o_222),
  .S0(dff_q_3)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_223),
  .I1(mux_o_224),
  .S0(dff_q_3)
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_225),
  .I1(mux_o_226),
  .S0(dff_q_3)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_227),
  .I1(mux_o_228),
  .S0(dff_q_3)
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(mux_o_229),
  .I1(mux_o_230),
  .S0(dff_q_3)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(dff_q_3)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(dff_q_2)
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_2)
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(dff_q_2)
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(mux_o_239),
  .I1(mux_o_240),
  .S0(dff_q_2)
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(mux_o_241),
  .I1(mux_o_242),
  .S0(dff_q_1)
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(mux_o_243),
  .I1(mux_o_244),
  .S0(dff_q_1)
);
MUX2 mux_inst_247 (
  .O(dout[7]),
  .I0(mux_o_245),
  .I1(mux_o_246),
  .S0(dff_q_0)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(sp_inst_0_dout[8]),
  .I1(sp_inst_1_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(sp_inst_2_dout[8]),
  .I1(sp_inst_3_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(sp_inst_4_dout[8]),
  .I1(sp_inst_5_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_251 (
  .O(mux_o_251),
  .I0(sp_inst_6_dout[8]),
  .I1(sp_inst_7_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(sp_inst_8_dout[8]),
  .I1(sp_inst_9_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(sp_inst_10_dout[8]),
  .I1(sp_inst_11_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(sp_inst_12_dout[8]),
  .I1(sp_inst_13_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(sp_inst_14_dout[8]),
  .I1(sp_inst_15_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(sp_inst_16_dout[8]),
  .I1(sp_inst_17_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(sp_inst_18_dout[8]),
  .I1(sp_inst_19_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(sp_inst_20_dout[8]),
  .I1(sp_inst_21_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(sp_inst_22_dout[8]),
  .I1(sp_inst_23_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(sp_inst_24_dout[8]),
  .I1(sp_inst_25_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(sp_inst_26_dout[8]),
  .I1(sp_inst_27_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(sp_inst_28_dout[8]),
  .I1(sp_inst_29_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(sp_inst_30_dout[8]),
  .I1(sp_inst_31_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(mux_o_248),
  .I1(mux_o_249),
  .S0(dff_q_3)
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(mux_o_250),
  .I1(mux_o_251),
  .S0(dff_q_3)
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(mux_o_252),
  .I1(mux_o_253),
  .S0(dff_q_3)
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(mux_o_254),
  .I1(mux_o_255),
  .S0(dff_q_3)
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(mux_o_256),
  .I1(mux_o_257),
  .S0(dff_q_3)
);
MUX2 mux_inst_269 (
  .O(mux_o_269),
  .I0(mux_o_258),
  .I1(mux_o_259),
  .S0(dff_q_3)
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(mux_o_260),
  .I1(mux_o_261),
  .S0(dff_q_3)
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(mux_o_262),
  .I1(mux_o_263),
  .S0(dff_q_3)
);
MUX2 mux_inst_272 (
  .O(mux_o_272),
  .I0(mux_o_264),
  .I1(mux_o_265),
  .S0(dff_q_2)
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(mux_o_266),
  .I1(mux_o_267),
  .S0(dff_q_2)
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(mux_o_268),
  .I1(mux_o_269),
  .S0(dff_q_2)
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(dff_q_2)
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(mux_o_272),
  .I1(mux_o_273),
  .S0(dff_q_1)
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(mux_o_274),
  .I1(mux_o_275),
  .S0(dff_q_1)
);
MUX2 mux_inst_278 (
  .O(dout[8]),
  .I0(mux_o_276),
  .I1(mux_o_277),
  .S0(dff_q_0)
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(sp_inst_0_dout[9]),
  .I1(sp_inst_1_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(sp_inst_2_dout[9]),
  .I1(sp_inst_3_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(sp_inst_4_dout[9]),
  .I1(sp_inst_5_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(sp_inst_6_dout[9]),
  .I1(sp_inst_7_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(sp_inst_8_dout[9]),
  .I1(sp_inst_9_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_284 (
  .O(mux_o_284),
  .I0(sp_inst_10_dout[9]),
  .I1(sp_inst_11_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(sp_inst_12_dout[9]),
  .I1(sp_inst_13_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(sp_inst_14_dout[9]),
  .I1(sp_inst_15_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(sp_inst_16_dout[9]),
  .I1(sp_inst_17_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(sp_inst_18_dout[9]),
  .I1(sp_inst_19_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(sp_inst_20_dout[9]),
  .I1(sp_inst_21_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(sp_inst_22_dout[9]),
  .I1(sp_inst_23_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(sp_inst_24_dout[9]),
  .I1(sp_inst_25_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(sp_inst_26_dout[9]),
  .I1(sp_inst_27_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(sp_inst_28_dout[9]),
  .I1(sp_inst_29_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(sp_inst_30_dout[9]),
  .I1(sp_inst_31_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(mux_o_279),
  .I1(mux_o_280),
  .S0(dff_q_3)
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(mux_o_281),
  .I1(mux_o_282),
  .S0(dff_q_3)
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(mux_o_283),
  .I1(mux_o_284),
  .S0(dff_q_3)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(mux_o_285),
  .I1(mux_o_286),
  .S0(dff_q_3)
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(mux_o_287),
  .I1(mux_o_288),
  .S0(dff_q_3)
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(mux_o_289),
  .I1(mux_o_290),
  .S0(dff_q_3)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(mux_o_291),
  .I1(mux_o_292),
  .S0(dff_q_3)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(mux_o_293),
  .I1(mux_o_294),
  .S0(dff_q_3)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(mux_o_295),
  .I1(mux_o_296),
  .S0(dff_q_2)
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(mux_o_297),
  .I1(mux_o_298),
  .S0(dff_q_2)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(mux_o_299),
  .I1(mux_o_300),
  .S0(dff_q_2)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(mux_o_301),
  .I1(mux_o_302),
  .S0(dff_q_2)
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(mux_o_303),
  .I1(mux_o_304),
  .S0(dff_q_1)
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(mux_o_305),
  .I1(mux_o_306),
  .S0(dff_q_1)
);
MUX2 mux_inst_309 (
  .O(dout[9]),
  .I0(mux_o_307),
  .I1(mux_o_308),
  .S0(dff_q_0)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(sp_inst_0_dout[10]),
  .I1(sp_inst_1_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(sp_inst_2_dout[10]),
  .I1(sp_inst_3_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(sp_inst_4_dout[10]),
  .I1(sp_inst_5_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(sp_inst_6_dout[10]),
  .I1(sp_inst_7_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_314 (
  .O(mux_o_314),
  .I0(sp_inst_8_dout[10]),
  .I1(sp_inst_9_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(sp_inst_10_dout[10]),
  .I1(sp_inst_11_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(sp_inst_12_dout[10]),
  .I1(sp_inst_13_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(sp_inst_14_dout[10]),
  .I1(sp_inst_15_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(sp_inst_16_dout[10]),
  .I1(sp_inst_17_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(sp_inst_18_dout[10]),
  .I1(sp_inst_19_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(sp_inst_20_dout[10]),
  .I1(sp_inst_21_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(sp_inst_22_dout[10]),
  .I1(sp_inst_23_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(sp_inst_24_dout[10]),
  .I1(sp_inst_25_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(sp_inst_26_dout[10]),
  .I1(sp_inst_27_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(sp_inst_28_dout[10]),
  .I1(sp_inst_29_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(sp_inst_30_dout[10]),
  .I1(sp_inst_31_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(dff_q_3)
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(dff_q_3)
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(mux_o_314),
  .I1(mux_o_315),
  .S0(dff_q_3)
);
MUX2 mux_inst_329 (
  .O(mux_o_329),
  .I0(mux_o_316),
  .I1(mux_o_317),
  .S0(dff_q_3)
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(mux_o_318),
  .I1(mux_o_319),
  .S0(dff_q_3)
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(mux_o_320),
  .I1(mux_o_321),
  .S0(dff_q_3)
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(mux_o_322),
  .I1(mux_o_323),
  .S0(dff_q_3)
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(mux_o_324),
  .I1(mux_o_325),
  .S0(dff_q_3)
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(mux_o_326),
  .I1(mux_o_327),
  .S0(dff_q_2)
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(mux_o_328),
  .I1(mux_o_329),
  .S0(dff_q_2)
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(mux_o_330),
  .I1(mux_o_331),
  .S0(dff_q_2)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(mux_o_332),
  .I1(mux_o_333),
  .S0(dff_q_2)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(mux_o_334),
  .I1(mux_o_335),
  .S0(dff_q_1)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(mux_o_336),
  .I1(mux_o_337),
  .S0(dff_q_1)
);
MUX2 mux_inst_340 (
  .O(dout[10]),
  .I0(mux_o_338),
  .I1(mux_o_339),
  .S0(dff_q_0)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(sp_inst_0_dout[11]),
  .I1(sp_inst_1_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(sp_inst_2_dout[11]),
  .I1(sp_inst_3_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(sp_inst_4_dout[11]),
  .I1(sp_inst_5_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(sp_inst_6_dout[11]),
  .I1(sp_inst_7_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(sp_inst_8_dout[11]),
  .I1(sp_inst_9_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(sp_inst_10_dout[11]),
  .I1(sp_inst_11_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(sp_inst_12_dout[11]),
  .I1(sp_inst_13_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(sp_inst_14_dout[11]),
  .I1(sp_inst_15_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_349 (
  .O(mux_o_349),
  .I0(sp_inst_16_dout[11]),
  .I1(sp_inst_17_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(sp_inst_18_dout[11]),
  .I1(sp_inst_19_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(sp_inst_20_dout[11]),
  .I1(sp_inst_21_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(sp_inst_22_dout[11]),
  .I1(sp_inst_23_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(sp_inst_24_dout[11]),
  .I1(sp_inst_25_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(sp_inst_26_dout[11]),
  .I1(sp_inst_27_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(sp_inst_28_dout[11]),
  .I1(sp_inst_29_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_356 (
  .O(mux_o_356),
  .I0(sp_inst_30_dout[11]),
  .I1(sp_inst_31_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_341),
  .I1(mux_o_342),
  .S0(dff_q_3)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_343),
  .I1(mux_o_344),
  .S0(dff_q_3)
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(mux_o_345),
  .I1(mux_o_346),
  .S0(dff_q_3)
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(dff_q_3)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_349),
  .I1(mux_o_350),
  .S0(dff_q_3)
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(mux_o_351),
  .I1(mux_o_352),
  .S0(dff_q_3)
);
MUX2 mux_inst_363 (
  .O(mux_o_363),
  .I0(mux_o_353),
  .I1(mux_o_354),
  .S0(dff_q_3)
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(mux_o_355),
  .I1(mux_o_356),
  .S0(dff_q_3)
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(dff_q_2)
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(mux_o_359),
  .I1(mux_o_360),
  .S0(dff_q_2)
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(mux_o_361),
  .I1(mux_o_362),
  .S0(dff_q_2)
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(mux_o_363),
  .I1(mux_o_364),
  .S0(dff_q_2)
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(mux_o_365),
  .I1(mux_o_366),
  .S0(dff_q_1)
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(mux_o_367),
  .I1(mux_o_368),
  .S0(dff_q_1)
);
MUX2 mux_inst_371 (
  .O(dout[11]),
  .I0(mux_o_369),
  .I1(mux_o_370),
  .S0(dff_q_0)
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(sp_inst_0_dout[12]),
  .I1(sp_inst_1_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(sp_inst_2_dout[12]),
  .I1(sp_inst_3_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_374 (
  .O(mux_o_374),
  .I0(sp_inst_4_dout[12]),
  .I1(sp_inst_5_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(sp_inst_6_dout[12]),
  .I1(sp_inst_7_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(sp_inst_8_dout[12]),
  .I1(sp_inst_9_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_377 (
  .O(mux_o_377),
  .I0(sp_inst_10_dout[12]),
  .I1(sp_inst_11_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_378 (
  .O(mux_o_378),
  .I0(sp_inst_12_dout[12]),
  .I1(sp_inst_13_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_379 (
  .O(mux_o_379),
  .I0(sp_inst_14_dout[12]),
  .I1(sp_inst_15_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_380 (
  .O(mux_o_380),
  .I0(sp_inst_16_dout[12]),
  .I1(sp_inst_17_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_381 (
  .O(mux_o_381),
  .I0(sp_inst_18_dout[12]),
  .I1(sp_inst_19_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_382 (
  .O(mux_o_382),
  .I0(sp_inst_20_dout[12]),
  .I1(sp_inst_21_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_383 (
  .O(mux_o_383),
  .I0(sp_inst_22_dout[12]),
  .I1(sp_inst_23_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_384 (
  .O(mux_o_384),
  .I0(sp_inst_24_dout[12]),
  .I1(sp_inst_25_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(sp_inst_26_dout[12]),
  .I1(sp_inst_27_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_386 (
  .O(mux_o_386),
  .I0(sp_inst_28_dout[12]),
  .I1(sp_inst_29_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_387 (
  .O(mux_o_387),
  .I0(sp_inst_30_dout[12]),
  .I1(sp_inst_31_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(mux_o_372),
  .I1(mux_o_373),
  .S0(dff_q_3)
);
MUX2 mux_inst_389 (
  .O(mux_o_389),
  .I0(mux_o_374),
  .I1(mux_o_375),
  .S0(dff_q_3)
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(mux_o_376),
  .I1(mux_o_377),
  .S0(dff_q_3)
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(mux_o_378),
  .I1(mux_o_379),
  .S0(dff_q_3)
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(mux_o_380),
  .I1(mux_o_381),
  .S0(dff_q_3)
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(mux_o_382),
  .I1(mux_o_383),
  .S0(dff_q_3)
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(mux_o_384),
  .I1(mux_o_385),
  .S0(dff_q_3)
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(mux_o_386),
  .I1(mux_o_387),
  .S0(dff_q_3)
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(mux_o_388),
  .I1(mux_o_389),
  .S0(dff_q_2)
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(mux_o_390),
  .I1(mux_o_391),
  .S0(dff_q_2)
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(mux_o_392),
  .I1(mux_o_393),
  .S0(dff_q_2)
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(mux_o_394),
  .I1(mux_o_395),
  .S0(dff_q_2)
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(mux_o_396),
  .I1(mux_o_397),
  .S0(dff_q_1)
);
MUX2 mux_inst_401 (
  .O(mux_o_401),
  .I0(mux_o_398),
  .I1(mux_o_399),
  .S0(dff_q_1)
);
MUX2 mux_inst_402 (
  .O(dout[12]),
  .I0(mux_o_400),
  .I1(mux_o_401),
  .S0(dff_q_0)
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(sp_inst_0_dout[13]),
  .I1(sp_inst_1_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_404 (
  .O(mux_o_404),
  .I0(sp_inst_2_dout[13]),
  .I1(sp_inst_3_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(sp_inst_4_dout[13]),
  .I1(sp_inst_5_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(sp_inst_6_dout[13]),
  .I1(sp_inst_7_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(sp_inst_8_dout[13]),
  .I1(sp_inst_9_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_408 (
  .O(mux_o_408),
  .I0(sp_inst_10_dout[13]),
  .I1(sp_inst_11_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(sp_inst_12_dout[13]),
  .I1(sp_inst_13_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(sp_inst_14_dout[13]),
  .I1(sp_inst_15_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(sp_inst_16_dout[13]),
  .I1(sp_inst_17_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_412 (
  .O(mux_o_412),
  .I0(sp_inst_18_dout[13]),
  .I1(sp_inst_19_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(sp_inst_20_dout[13]),
  .I1(sp_inst_21_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(sp_inst_22_dout[13]),
  .I1(sp_inst_23_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_415 (
  .O(mux_o_415),
  .I0(sp_inst_24_dout[13]),
  .I1(sp_inst_25_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_416 (
  .O(mux_o_416),
  .I0(sp_inst_26_dout[13]),
  .I1(sp_inst_27_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_417 (
  .O(mux_o_417),
  .I0(sp_inst_28_dout[13]),
  .I1(sp_inst_29_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_418 (
  .O(mux_o_418),
  .I0(sp_inst_30_dout[13]),
  .I1(sp_inst_31_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_419 (
  .O(mux_o_419),
  .I0(mux_o_403),
  .I1(mux_o_404),
  .S0(dff_q_3)
);
MUX2 mux_inst_420 (
  .O(mux_o_420),
  .I0(mux_o_405),
  .I1(mux_o_406),
  .S0(dff_q_3)
);
MUX2 mux_inst_421 (
  .O(mux_o_421),
  .I0(mux_o_407),
  .I1(mux_o_408),
  .S0(dff_q_3)
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(mux_o_409),
  .I1(mux_o_410),
  .S0(dff_q_3)
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(mux_o_411),
  .I1(mux_o_412),
  .S0(dff_q_3)
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(mux_o_413),
  .I1(mux_o_414),
  .S0(dff_q_3)
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(mux_o_415),
  .I1(mux_o_416),
  .S0(dff_q_3)
);
MUX2 mux_inst_426 (
  .O(mux_o_426),
  .I0(mux_o_417),
  .I1(mux_o_418),
  .S0(dff_q_3)
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(mux_o_419),
  .I1(mux_o_420),
  .S0(dff_q_2)
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(mux_o_421),
  .I1(mux_o_422),
  .S0(dff_q_2)
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(mux_o_423),
  .I1(mux_o_424),
  .S0(dff_q_2)
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(mux_o_425),
  .I1(mux_o_426),
  .S0(dff_q_2)
);
MUX2 mux_inst_431 (
  .O(mux_o_431),
  .I0(mux_o_427),
  .I1(mux_o_428),
  .S0(dff_q_1)
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(mux_o_429),
  .I1(mux_o_430),
  .S0(dff_q_1)
);
MUX2 mux_inst_433 (
  .O(dout[13]),
  .I0(mux_o_431),
  .I1(mux_o_432),
  .S0(dff_q_0)
);
MUX2 mux_inst_434 (
  .O(mux_o_434),
  .I0(sp_inst_0_dout[14]),
  .I1(sp_inst_1_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(sp_inst_2_dout[14]),
  .I1(sp_inst_3_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(sp_inst_4_dout[14]),
  .I1(sp_inst_5_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(sp_inst_6_dout[14]),
  .I1(sp_inst_7_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(sp_inst_8_dout[14]),
  .I1(sp_inst_9_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(sp_inst_10_dout[14]),
  .I1(sp_inst_11_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_440 (
  .O(mux_o_440),
  .I0(sp_inst_12_dout[14]),
  .I1(sp_inst_13_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(sp_inst_14_dout[14]),
  .I1(sp_inst_15_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(sp_inst_16_dout[14]),
  .I1(sp_inst_17_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(sp_inst_18_dout[14]),
  .I1(sp_inst_19_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(sp_inst_20_dout[14]),
  .I1(sp_inst_21_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(sp_inst_22_dout[14]),
  .I1(sp_inst_23_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(sp_inst_24_dout[14]),
  .I1(sp_inst_25_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(sp_inst_26_dout[14]),
  .I1(sp_inst_27_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(sp_inst_28_dout[14]),
  .I1(sp_inst_29_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_449 (
  .O(mux_o_449),
  .I0(sp_inst_30_dout[14]),
  .I1(sp_inst_31_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(mux_o_434),
  .I1(mux_o_435),
  .S0(dff_q_3)
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(mux_o_436),
  .I1(mux_o_437),
  .S0(dff_q_3)
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(mux_o_438),
  .I1(mux_o_439),
  .S0(dff_q_3)
);
MUX2 mux_inst_453 (
  .O(mux_o_453),
  .I0(mux_o_440),
  .I1(mux_o_441),
  .S0(dff_q_3)
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(mux_o_442),
  .I1(mux_o_443),
  .S0(dff_q_3)
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(mux_o_444),
  .I1(mux_o_445),
  .S0(dff_q_3)
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(mux_o_446),
  .I1(mux_o_447),
  .S0(dff_q_3)
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(mux_o_448),
  .I1(mux_o_449),
  .S0(dff_q_3)
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(mux_o_450),
  .I1(mux_o_451),
  .S0(dff_q_2)
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(mux_o_452),
  .I1(mux_o_453),
  .S0(dff_q_2)
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(mux_o_454),
  .I1(mux_o_455),
  .S0(dff_q_2)
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(mux_o_456),
  .I1(mux_o_457),
  .S0(dff_q_2)
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(mux_o_458),
  .I1(mux_o_459),
  .S0(dff_q_1)
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(mux_o_460),
  .I1(mux_o_461),
  .S0(dff_q_1)
);
MUX2 mux_inst_464 (
  .O(dout[14]),
  .I0(mux_o_462),
  .I1(mux_o_463),
  .S0(dff_q_0)
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(sp_inst_0_dout[15]),
  .I1(sp_inst_1_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(sp_inst_2_dout[15]),
  .I1(sp_inst_3_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_467 (
  .O(mux_o_467),
  .I0(sp_inst_4_dout[15]),
  .I1(sp_inst_5_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_468 (
  .O(mux_o_468),
  .I0(sp_inst_6_dout[15]),
  .I1(sp_inst_7_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_469 (
  .O(mux_o_469),
  .I0(sp_inst_8_dout[15]),
  .I1(sp_inst_9_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_470 (
  .O(mux_o_470),
  .I0(sp_inst_10_dout[15]),
  .I1(sp_inst_11_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_471 (
  .O(mux_o_471),
  .I0(sp_inst_12_dout[15]),
  .I1(sp_inst_13_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(sp_inst_14_dout[15]),
  .I1(sp_inst_15_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_473 (
  .O(mux_o_473),
  .I0(sp_inst_16_dout[15]),
  .I1(sp_inst_17_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_474 (
  .O(mux_o_474),
  .I0(sp_inst_18_dout[15]),
  .I1(sp_inst_19_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_475 (
  .O(mux_o_475),
  .I0(sp_inst_20_dout[15]),
  .I1(sp_inst_21_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_476 (
  .O(mux_o_476),
  .I0(sp_inst_22_dout[15]),
  .I1(sp_inst_23_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_477 (
  .O(mux_o_477),
  .I0(sp_inst_24_dout[15]),
  .I1(sp_inst_25_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_478 (
  .O(mux_o_478),
  .I0(sp_inst_26_dout[15]),
  .I1(sp_inst_27_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_479 (
  .O(mux_o_479),
  .I0(sp_inst_28_dout[15]),
  .I1(sp_inst_29_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_480 (
  .O(mux_o_480),
  .I0(sp_inst_30_dout[15]),
  .I1(sp_inst_31_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_481 (
  .O(mux_o_481),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(dff_q_3)
);
MUX2 mux_inst_482 (
  .O(mux_o_482),
  .I0(mux_o_467),
  .I1(mux_o_468),
  .S0(dff_q_3)
);
MUX2 mux_inst_483 (
  .O(mux_o_483),
  .I0(mux_o_469),
  .I1(mux_o_470),
  .S0(dff_q_3)
);
MUX2 mux_inst_484 (
  .O(mux_o_484),
  .I0(mux_o_471),
  .I1(mux_o_472),
  .S0(dff_q_3)
);
MUX2 mux_inst_485 (
  .O(mux_o_485),
  .I0(mux_o_473),
  .I1(mux_o_474),
  .S0(dff_q_3)
);
MUX2 mux_inst_486 (
  .O(mux_o_486),
  .I0(mux_o_475),
  .I1(mux_o_476),
  .S0(dff_q_3)
);
MUX2 mux_inst_487 (
  .O(mux_o_487),
  .I0(mux_o_477),
  .I1(mux_o_478),
  .S0(dff_q_3)
);
MUX2 mux_inst_488 (
  .O(mux_o_488),
  .I0(mux_o_479),
  .I1(mux_o_480),
  .S0(dff_q_3)
);
MUX2 mux_inst_489 (
  .O(mux_o_489),
  .I0(mux_o_481),
  .I1(mux_o_482),
  .S0(dff_q_2)
);
MUX2 mux_inst_490 (
  .O(mux_o_490),
  .I0(mux_o_483),
  .I1(mux_o_484),
  .S0(dff_q_2)
);
MUX2 mux_inst_491 (
  .O(mux_o_491),
  .I0(mux_o_485),
  .I1(mux_o_486),
  .S0(dff_q_2)
);
MUX2 mux_inst_492 (
  .O(mux_o_492),
  .I0(mux_o_487),
  .I1(mux_o_488),
  .S0(dff_q_2)
);
MUX2 mux_inst_493 (
  .O(mux_o_493),
  .I0(mux_o_489),
  .I1(mux_o_490),
  .S0(dff_q_1)
);
MUX2 mux_inst_494 (
  .O(mux_o_494),
  .I0(mux_o_491),
  .I1(mux_o_492),
  .S0(dff_q_1)
);
MUX2 mux_inst_495 (
  .O(dout[15]),
  .I0(mux_o_493),
  .I1(mux_o_494),
  .S0(dff_q_0)
);
MUX2 mux_inst_496 (
  .O(mux_o_496),
  .I0(sp_inst_32_dout[16]),
  .I1(sp_inst_33_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_497 (
  .O(mux_o_497),
  .I0(sp_inst_34_dout[16]),
  .I1(sp_inst_35_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_498 (
  .O(mux_o_498),
  .I0(sp_inst_36_dout[16]),
  .I1(sp_inst_37_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_499 (
  .O(mux_o_499),
  .I0(sp_inst_38_dout[16]),
  .I1(sp_inst_39_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_500 (
  .O(mux_o_500),
  .I0(sp_inst_40_dout[16]),
  .I1(sp_inst_41_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_501 (
  .O(mux_o_501),
  .I0(sp_inst_42_dout[16]),
  .I1(sp_inst_43_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_502 (
  .O(mux_o_502),
  .I0(sp_inst_44_dout[16]),
  .I1(sp_inst_45_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_503 (
  .O(mux_o_503),
  .I0(sp_inst_46_dout[16]),
  .I1(sp_inst_47_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_504 (
  .O(mux_o_504),
  .I0(sp_inst_48_dout[16]),
  .I1(sp_inst_49_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_505 (
  .O(mux_o_505),
  .I0(sp_inst_50_dout[16]),
  .I1(sp_inst_51_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_506 (
  .O(mux_o_506),
  .I0(sp_inst_52_dout[16]),
  .I1(sp_inst_53_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_507 (
  .O(mux_o_507),
  .I0(sp_inst_54_dout[16]),
  .I1(sp_inst_55_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_508 (
  .O(mux_o_508),
  .I0(sp_inst_56_dout[16]),
  .I1(sp_inst_57_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_509 (
  .O(mux_o_509),
  .I0(sp_inst_58_dout[16]),
  .I1(sp_inst_59_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_510 (
  .O(mux_o_510),
  .I0(sp_inst_60_dout[16]),
  .I1(sp_inst_61_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_511 (
  .O(mux_o_511),
  .I0(sp_inst_62_dout[16]),
  .I1(sp_inst_63_dout[16]),
  .S0(dff_q_4)
);
MUX2 mux_inst_512 (
  .O(mux_o_512),
  .I0(mux_o_496),
  .I1(mux_o_497),
  .S0(dff_q_3)
);
MUX2 mux_inst_513 (
  .O(mux_o_513),
  .I0(mux_o_498),
  .I1(mux_o_499),
  .S0(dff_q_3)
);
MUX2 mux_inst_514 (
  .O(mux_o_514),
  .I0(mux_o_500),
  .I1(mux_o_501),
  .S0(dff_q_3)
);
MUX2 mux_inst_515 (
  .O(mux_o_515),
  .I0(mux_o_502),
  .I1(mux_o_503),
  .S0(dff_q_3)
);
MUX2 mux_inst_516 (
  .O(mux_o_516),
  .I0(mux_o_504),
  .I1(mux_o_505),
  .S0(dff_q_3)
);
MUX2 mux_inst_517 (
  .O(mux_o_517),
  .I0(mux_o_506),
  .I1(mux_o_507),
  .S0(dff_q_3)
);
MUX2 mux_inst_518 (
  .O(mux_o_518),
  .I0(mux_o_508),
  .I1(mux_o_509),
  .S0(dff_q_3)
);
MUX2 mux_inst_519 (
  .O(mux_o_519),
  .I0(mux_o_510),
  .I1(mux_o_511),
  .S0(dff_q_3)
);
MUX2 mux_inst_520 (
  .O(mux_o_520),
  .I0(mux_o_512),
  .I1(mux_o_513),
  .S0(dff_q_2)
);
MUX2 mux_inst_521 (
  .O(mux_o_521),
  .I0(mux_o_514),
  .I1(mux_o_515),
  .S0(dff_q_2)
);
MUX2 mux_inst_522 (
  .O(mux_o_522),
  .I0(mux_o_516),
  .I1(mux_o_517),
  .S0(dff_q_2)
);
MUX2 mux_inst_523 (
  .O(mux_o_523),
  .I0(mux_o_518),
  .I1(mux_o_519),
  .S0(dff_q_2)
);
MUX2 mux_inst_524 (
  .O(mux_o_524),
  .I0(mux_o_520),
  .I1(mux_o_521),
  .S0(dff_q_1)
);
MUX2 mux_inst_525 (
  .O(mux_o_525),
  .I0(mux_o_522),
  .I1(mux_o_523),
  .S0(dff_q_1)
);
MUX2 mux_inst_526 (
  .O(dout[16]),
  .I0(mux_o_524),
  .I1(mux_o_525),
  .S0(dff_q_0)
);
MUX2 mux_inst_527 (
  .O(mux_o_527),
  .I0(sp_inst_32_dout[17]),
  .I1(sp_inst_33_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_528 (
  .O(mux_o_528),
  .I0(sp_inst_34_dout[17]),
  .I1(sp_inst_35_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_529 (
  .O(mux_o_529),
  .I0(sp_inst_36_dout[17]),
  .I1(sp_inst_37_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_530 (
  .O(mux_o_530),
  .I0(sp_inst_38_dout[17]),
  .I1(sp_inst_39_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_531 (
  .O(mux_o_531),
  .I0(sp_inst_40_dout[17]),
  .I1(sp_inst_41_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_532 (
  .O(mux_o_532),
  .I0(sp_inst_42_dout[17]),
  .I1(sp_inst_43_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_533 (
  .O(mux_o_533),
  .I0(sp_inst_44_dout[17]),
  .I1(sp_inst_45_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_534 (
  .O(mux_o_534),
  .I0(sp_inst_46_dout[17]),
  .I1(sp_inst_47_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_535 (
  .O(mux_o_535),
  .I0(sp_inst_48_dout[17]),
  .I1(sp_inst_49_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_536 (
  .O(mux_o_536),
  .I0(sp_inst_50_dout[17]),
  .I1(sp_inst_51_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_537 (
  .O(mux_o_537),
  .I0(sp_inst_52_dout[17]),
  .I1(sp_inst_53_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_538 (
  .O(mux_o_538),
  .I0(sp_inst_54_dout[17]),
  .I1(sp_inst_55_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_539 (
  .O(mux_o_539),
  .I0(sp_inst_56_dout[17]),
  .I1(sp_inst_57_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_540 (
  .O(mux_o_540),
  .I0(sp_inst_58_dout[17]),
  .I1(sp_inst_59_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_541 (
  .O(mux_o_541),
  .I0(sp_inst_60_dout[17]),
  .I1(sp_inst_61_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_542 (
  .O(mux_o_542),
  .I0(sp_inst_62_dout[17]),
  .I1(sp_inst_63_dout[17]),
  .S0(dff_q_4)
);
MUX2 mux_inst_543 (
  .O(mux_o_543),
  .I0(mux_o_527),
  .I1(mux_o_528),
  .S0(dff_q_3)
);
MUX2 mux_inst_544 (
  .O(mux_o_544),
  .I0(mux_o_529),
  .I1(mux_o_530),
  .S0(dff_q_3)
);
MUX2 mux_inst_545 (
  .O(mux_o_545),
  .I0(mux_o_531),
  .I1(mux_o_532),
  .S0(dff_q_3)
);
MUX2 mux_inst_546 (
  .O(mux_o_546),
  .I0(mux_o_533),
  .I1(mux_o_534),
  .S0(dff_q_3)
);
MUX2 mux_inst_547 (
  .O(mux_o_547),
  .I0(mux_o_535),
  .I1(mux_o_536),
  .S0(dff_q_3)
);
MUX2 mux_inst_548 (
  .O(mux_o_548),
  .I0(mux_o_537),
  .I1(mux_o_538),
  .S0(dff_q_3)
);
MUX2 mux_inst_549 (
  .O(mux_o_549),
  .I0(mux_o_539),
  .I1(mux_o_540),
  .S0(dff_q_3)
);
MUX2 mux_inst_550 (
  .O(mux_o_550),
  .I0(mux_o_541),
  .I1(mux_o_542),
  .S0(dff_q_3)
);
MUX2 mux_inst_551 (
  .O(mux_o_551),
  .I0(mux_o_543),
  .I1(mux_o_544),
  .S0(dff_q_2)
);
MUX2 mux_inst_552 (
  .O(mux_o_552),
  .I0(mux_o_545),
  .I1(mux_o_546),
  .S0(dff_q_2)
);
MUX2 mux_inst_553 (
  .O(mux_o_553),
  .I0(mux_o_547),
  .I1(mux_o_548),
  .S0(dff_q_2)
);
MUX2 mux_inst_554 (
  .O(mux_o_554),
  .I0(mux_o_549),
  .I1(mux_o_550),
  .S0(dff_q_2)
);
MUX2 mux_inst_555 (
  .O(mux_o_555),
  .I0(mux_o_551),
  .I1(mux_o_552),
  .S0(dff_q_1)
);
MUX2 mux_inst_556 (
  .O(mux_o_556),
  .I0(mux_o_553),
  .I1(mux_o_554),
  .S0(dff_q_1)
);
MUX2 mux_inst_557 (
  .O(dout[17]),
  .I0(mux_o_555),
  .I1(mux_o_556),
  .S0(dff_q_0)
);
MUX2 mux_inst_558 (
  .O(mux_o_558),
  .I0(sp_inst_32_dout[18]),
  .I1(sp_inst_33_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_559 (
  .O(mux_o_559),
  .I0(sp_inst_34_dout[18]),
  .I1(sp_inst_35_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_560 (
  .O(mux_o_560),
  .I0(sp_inst_36_dout[18]),
  .I1(sp_inst_37_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_561 (
  .O(mux_o_561),
  .I0(sp_inst_38_dout[18]),
  .I1(sp_inst_39_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_562 (
  .O(mux_o_562),
  .I0(sp_inst_40_dout[18]),
  .I1(sp_inst_41_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_563 (
  .O(mux_o_563),
  .I0(sp_inst_42_dout[18]),
  .I1(sp_inst_43_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_564 (
  .O(mux_o_564),
  .I0(sp_inst_44_dout[18]),
  .I1(sp_inst_45_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_565 (
  .O(mux_o_565),
  .I0(sp_inst_46_dout[18]),
  .I1(sp_inst_47_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_566 (
  .O(mux_o_566),
  .I0(sp_inst_48_dout[18]),
  .I1(sp_inst_49_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_567 (
  .O(mux_o_567),
  .I0(sp_inst_50_dout[18]),
  .I1(sp_inst_51_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_568 (
  .O(mux_o_568),
  .I0(sp_inst_52_dout[18]),
  .I1(sp_inst_53_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_569 (
  .O(mux_o_569),
  .I0(sp_inst_54_dout[18]),
  .I1(sp_inst_55_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_570 (
  .O(mux_o_570),
  .I0(sp_inst_56_dout[18]),
  .I1(sp_inst_57_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_571 (
  .O(mux_o_571),
  .I0(sp_inst_58_dout[18]),
  .I1(sp_inst_59_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_572 (
  .O(mux_o_572),
  .I0(sp_inst_60_dout[18]),
  .I1(sp_inst_61_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_573 (
  .O(mux_o_573),
  .I0(sp_inst_62_dout[18]),
  .I1(sp_inst_63_dout[18]),
  .S0(dff_q_4)
);
MUX2 mux_inst_574 (
  .O(mux_o_574),
  .I0(mux_o_558),
  .I1(mux_o_559),
  .S0(dff_q_3)
);
MUX2 mux_inst_575 (
  .O(mux_o_575),
  .I0(mux_o_560),
  .I1(mux_o_561),
  .S0(dff_q_3)
);
MUX2 mux_inst_576 (
  .O(mux_o_576),
  .I0(mux_o_562),
  .I1(mux_o_563),
  .S0(dff_q_3)
);
MUX2 mux_inst_577 (
  .O(mux_o_577),
  .I0(mux_o_564),
  .I1(mux_o_565),
  .S0(dff_q_3)
);
MUX2 mux_inst_578 (
  .O(mux_o_578),
  .I0(mux_o_566),
  .I1(mux_o_567),
  .S0(dff_q_3)
);
MUX2 mux_inst_579 (
  .O(mux_o_579),
  .I0(mux_o_568),
  .I1(mux_o_569),
  .S0(dff_q_3)
);
MUX2 mux_inst_580 (
  .O(mux_o_580),
  .I0(mux_o_570),
  .I1(mux_o_571),
  .S0(dff_q_3)
);
MUX2 mux_inst_581 (
  .O(mux_o_581),
  .I0(mux_o_572),
  .I1(mux_o_573),
  .S0(dff_q_3)
);
MUX2 mux_inst_582 (
  .O(mux_o_582),
  .I0(mux_o_574),
  .I1(mux_o_575),
  .S0(dff_q_2)
);
MUX2 mux_inst_583 (
  .O(mux_o_583),
  .I0(mux_o_576),
  .I1(mux_o_577),
  .S0(dff_q_2)
);
MUX2 mux_inst_584 (
  .O(mux_o_584),
  .I0(mux_o_578),
  .I1(mux_o_579),
  .S0(dff_q_2)
);
MUX2 mux_inst_585 (
  .O(mux_o_585),
  .I0(mux_o_580),
  .I1(mux_o_581),
  .S0(dff_q_2)
);
MUX2 mux_inst_586 (
  .O(mux_o_586),
  .I0(mux_o_582),
  .I1(mux_o_583),
  .S0(dff_q_1)
);
MUX2 mux_inst_587 (
  .O(mux_o_587),
  .I0(mux_o_584),
  .I1(mux_o_585),
  .S0(dff_q_1)
);
MUX2 mux_inst_588 (
  .O(dout[18]),
  .I0(mux_o_586),
  .I1(mux_o_587),
  .S0(dff_q_0)
);
MUX2 mux_inst_589 (
  .O(mux_o_589),
  .I0(sp_inst_32_dout[19]),
  .I1(sp_inst_33_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_590 (
  .O(mux_o_590),
  .I0(sp_inst_34_dout[19]),
  .I1(sp_inst_35_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_591 (
  .O(mux_o_591),
  .I0(sp_inst_36_dout[19]),
  .I1(sp_inst_37_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_592 (
  .O(mux_o_592),
  .I0(sp_inst_38_dout[19]),
  .I1(sp_inst_39_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_593 (
  .O(mux_o_593),
  .I0(sp_inst_40_dout[19]),
  .I1(sp_inst_41_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_594 (
  .O(mux_o_594),
  .I0(sp_inst_42_dout[19]),
  .I1(sp_inst_43_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_595 (
  .O(mux_o_595),
  .I0(sp_inst_44_dout[19]),
  .I1(sp_inst_45_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_596 (
  .O(mux_o_596),
  .I0(sp_inst_46_dout[19]),
  .I1(sp_inst_47_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_597 (
  .O(mux_o_597),
  .I0(sp_inst_48_dout[19]),
  .I1(sp_inst_49_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_598 (
  .O(mux_o_598),
  .I0(sp_inst_50_dout[19]),
  .I1(sp_inst_51_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_599 (
  .O(mux_o_599),
  .I0(sp_inst_52_dout[19]),
  .I1(sp_inst_53_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_600 (
  .O(mux_o_600),
  .I0(sp_inst_54_dout[19]),
  .I1(sp_inst_55_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_601 (
  .O(mux_o_601),
  .I0(sp_inst_56_dout[19]),
  .I1(sp_inst_57_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_602 (
  .O(mux_o_602),
  .I0(sp_inst_58_dout[19]),
  .I1(sp_inst_59_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_603 (
  .O(mux_o_603),
  .I0(sp_inst_60_dout[19]),
  .I1(sp_inst_61_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_604 (
  .O(mux_o_604),
  .I0(sp_inst_62_dout[19]),
  .I1(sp_inst_63_dout[19]),
  .S0(dff_q_4)
);
MUX2 mux_inst_605 (
  .O(mux_o_605),
  .I0(mux_o_589),
  .I1(mux_o_590),
  .S0(dff_q_3)
);
MUX2 mux_inst_606 (
  .O(mux_o_606),
  .I0(mux_o_591),
  .I1(mux_o_592),
  .S0(dff_q_3)
);
MUX2 mux_inst_607 (
  .O(mux_o_607),
  .I0(mux_o_593),
  .I1(mux_o_594),
  .S0(dff_q_3)
);
MUX2 mux_inst_608 (
  .O(mux_o_608),
  .I0(mux_o_595),
  .I1(mux_o_596),
  .S0(dff_q_3)
);
MUX2 mux_inst_609 (
  .O(mux_o_609),
  .I0(mux_o_597),
  .I1(mux_o_598),
  .S0(dff_q_3)
);
MUX2 mux_inst_610 (
  .O(mux_o_610),
  .I0(mux_o_599),
  .I1(mux_o_600),
  .S0(dff_q_3)
);
MUX2 mux_inst_611 (
  .O(mux_o_611),
  .I0(mux_o_601),
  .I1(mux_o_602),
  .S0(dff_q_3)
);
MUX2 mux_inst_612 (
  .O(mux_o_612),
  .I0(mux_o_603),
  .I1(mux_o_604),
  .S0(dff_q_3)
);
MUX2 mux_inst_613 (
  .O(mux_o_613),
  .I0(mux_o_605),
  .I1(mux_o_606),
  .S0(dff_q_2)
);
MUX2 mux_inst_614 (
  .O(mux_o_614),
  .I0(mux_o_607),
  .I1(mux_o_608),
  .S0(dff_q_2)
);
MUX2 mux_inst_615 (
  .O(mux_o_615),
  .I0(mux_o_609),
  .I1(mux_o_610),
  .S0(dff_q_2)
);
MUX2 mux_inst_616 (
  .O(mux_o_616),
  .I0(mux_o_611),
  .I1(mux_o_612),
  .S0(dff_q_2)
);
MUX2 mux_inst_617 (
  .O(mux_o_617),
  .I0(mux_o_613),
  .I1(mux_o_614),
  .S0(dff_q_1)
);
MUX2 mux_inst_618 (
  .O(mux_o_618),
  .I0(mux_o_615),
  .I1(mux_o_616),
  .S0(dff_q_1)
);
MUX2 mux_inst_619 (
  .O(dout[19]),
  .I0(mux_o_617),
  .I1(mux_o_618),
  .S0(dff_q_0)
);
MUX2 mux_inst_620 (
  .O(mux_o_620),
  .I0(sp_inst_32_dout[20]),
  .I1(sp_inst_33_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_621 (
  .O(mux_o_621),
  .I0(sp_inst_34_dout[20]),
  .I1(sp_inst_35_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_622 (
  .O(mux_o_622),
  .I0(sp_inst_36_dout[20]),
  .I1(sp_inst_37_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_623 (
  .O(mux_o_623),
  .I0(sp_inst_38_dout[20]),
  .I1(sp_inst_39_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_624 (
  .O(mux_o_624),
  .I0(sp_inst_40_dout[20]),
  .I1(sp_inst_41_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_625 (
  .O(mux_o_625),
  .I0(sp_inst_42_dout[20]),
  .I1(sp_inst_43_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_626 (
  .O(mux_o_626),
  .I0(sp_inst_44_dout[20]),
  .I1(sp_inst_45_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_627 (
  .O(mux_o_627),
  .I0(sp_inst_46_dout[20]),
  .I1(sp_inst_47_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_628 (
  .O(mux_o_628),
  .I0(sp_inst_48_dout[20]),
  .I1(sp_inst_49_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_629 (
  .O(mux_o_629),
  .I0(sp_inst_50_dout[20]),
  .I1(sp_inst_51_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_630 (
  .O(mux_o_630),
  .I0(sp_inst_52_dout[20]),
  .I1(sp_inst_53_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_631 (
  .O(mux_o_631),
  .I0(sp_inst_54_dout[20]),
  .I1(sp_inst_55_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_632 (
  .O(mux_o_632),
  .I0(sp_inst_56_dout[20]),
  .I1(sp_inst_57_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_633 (
  .O(mux_o_633),
  .I0(sp_inst_58_dout[20]),
  .I1(sp_inst_59_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_634 (
  .O(mux_o_634),
  .I0(sp_inst_60_dout[20]),
  .I1(sp_inst_61_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_635 (
  .O(mux_o_635),
  .I0(sp_inst_62_dout[20]),
  .I1(sp_inst_63_dout[20]),
  .S0(dff_q_4)
);
MUX2 mux_inst_636 (
  .O(mux_o_636),
  .I0(mux_o_620),
  .I1(mux_o_621),
  .S0(dff_q_3)
);
MUX2 mux_inst_637 (
  .O(mux_o_637),
  .I0(mux_o_622),
  .I1(mux_o_623),
  .S0(dff_q_3)
);
MUX2 mux_inst_638 (
  .O(mux_o_638),
  .I0(mux_o_624),
  .I1(mux_o_625),
  .S0(dff_q_3)
);
MUX2 mux_inst_639 (
  .O(mux_o_639),
  .I0(mux_o_626),
  .I1(mux_o_627),
  .S0(dff_q_3)
);
MUX2 mux_inst_640 (
  .O(mux_o_640),
  .I0(mux_o_628),
  .I1(mux_o_629),
  .S0(dff_q_3)
);
MUX2 mux_inst_641 (
  .O(mux_o_641),
  .I0(mux_o_630),
  .I1(mux_o_631),
  .S0(dff_q_3)
);
MUX2 mux_inst_642 (
  .O(mux_o_642),
  .I0(mux_o_632),
  .I1(mux_o_633),
  .S0(dff_q_3)
);
MUX2 mux_inst_643 (
  .O(mux_o_643),
  .I0(mux_o_634),
  .I1(mux_o_635),
  .S0(dff_q_3)
);
MUX2 mux_inst_644 (
  .O(mux_o_644),
  .I0(mux_o_636),
  .I1(mux_o_637),
  .S0(dff_q_2)
);
MUX2 mux_inst_645 (
  .O(mux_o_645),
  .I0(mux_o_638),
  .I1(mux_o_639),
  .S0(dff_q_2)
);
MUX2 mux_inst_646 (
  .O(mux_o_646),
  .I0(mux_o_640),
  .I1(mux_o_641),
  .S0(dff_q_2)
);
MUX2 mux_inst_647 (
  .O(mux_o_647),
  .I0(mux_o_642),
  .I1(mux_o_643),
  .S0(dff_q_2)
);
MUX2 mux_inst_648 (
  .O(mux_o_648),
  .I0(mux_o_644),
  .I1(mux_o_645),
  .S0(dff_q_1)
);
MUX2 mux_inst_649 (
  .O(mux_o_649),
  .I0(mux_o_646),
  .I1(mux_o_647),
  .S0(dff_q_1)
);
MUX2 mux_inst_650 (
  .O(dout[20]),
  .I0(mux_o_648),
  .I1(mux_o_649),
  .S0(dff_q_0)
);
MUX2 mux_inst_651 (
  .O(mux_o_651),
  .I0(sp_inst_32_dout[21]),
  .I1(sp_inst_33_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_652 (
  .O(mux_o_652),
  .I0(sp_inst_34_dout[21]),
  .I1(sp_inst_35_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_653 (
  .O(mux_o_653),
  .I0(sp_inst_36_dout[21]),
  .I1(sp_inst_37_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_654 (
  .O(mux_o_654),
  .I0(sp_inst_38_dout[21]),
  .I1(sp_inst_39_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_655 (
  .O(mux_o_655),
  .I0(sp_inst_40_dout[21]),
  .I1(sp_inst_41_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_656 (
  .O(mux_o_656),
  .I0(sp_inst_42_dout[21]),
  .I1(sp_inst_43_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_657 (
  .O(mux_o_657),
  .I0(sp_inst_44_dout[21]),
  .I1(sp_inst_45_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_658 (
  .O(mux_o_658),
  .I0(sp_inst_46_dout[21]),
  .I1(sp_inst_47_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_659 (
  .O(mux_o_659),
  .I0(sp_inst_48_dout[21]),
  .I1(sp_inst_49_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_660 (
  .O(mux_o_660),
  .I0(sp_inst_50_dout[21]),
  .I1(sp_inst_51_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_661 (
  .O(mux_o_661),
  .I0(sp_inst_52_dout[21]),
  .I1(sp_inst_53_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_662 (
  .O(mux_o_662),
  .I0(sp_inst_54_dout[21]),
  .I1(sp_inst_55_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_663 (
  .O(mux_o_663),
  .I0(sp_inst_56_dout[21]),
  .I1(sp_inst_57_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_664 (
  .O(mux_o_664),
  .I0(sp_inst_58_dout[21]),
  .I1(sp_inst_59_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_665 (
  .O(mux_o_665),
  .I0(sp_inst_60_dout[21]),
  .I1(sp_inst_61_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_666 (
  .O(mux_o_666),
  .I0(sp_inst_62_dout[21]),
  .I1(sp_inst_63_dout[21]),
  .S0(dff_q_4)
);
MUX2 mux_inst_667 (
  .O(mux_o_667),
  .I0(mux_o_651),
  .I1(mux_o_652),
  .S0(dff_q_3)
);
MUX2 mux_inst_668 (
  .O(mux_o_668),
  .I0(mux_o_653),
  .I1(mux_o_654),
  .S0(dff_q_3)
);
MUX2 mux_inst_669 (
  .O(mux_o_669),
  .I0(mux_o_655),
  .I1(mux_o_656),
  .S0(dff_q_3)
);
MUX2 mux_inst_670 (
  .O(mux_o_670),
  .I0(mux_o_657),
  .I1(mux_o_658),
  .S0(dff_q_3)
);
MUX2 mux_inst_671 (
  .O(mux_o_671),
  .I0(mux_o_659),
  .I1(mux_o_660),
  .S0(dff_q_3)
);
MUX2 mux_inst_672 (
  .O(mux_o_672),
  .I0(mux_o_661),
  .I1(mux_o_662),
  .S0(dff_q_3)
);
MUX2 mux_inst_673 (
  .O(mux_o_673),
  .I0(mux_o_663),
  .I1(mux_o_664),
  .S0(dff_q_3)
);
MUX2 mux_inst_674 (
  .O(mux_o_674),
  .I0(mux_o_665),
  .I1(mux_o_666),
  .S0(dff_q_3)
);
MUX2 mux_inst_675 (
  .O(mux_o_675),
  .I0(mux_o_667),
  .I1(mux_o_668),
  .S0(dff_q_2)
);
MUX2 mux_inst_676 (
  .O(mux_o_676),
  .I0(mux_o_669),
  .I1(mux_o_670),
  .S0(dff_q_2)
);
MUX2 mux_inst_677 (
  .O(mux_o_677),
  .I0(mux_o_671),
  .I1(mux_o_672),
  .S0(dff_q_2)
);
MUX2 mux_inst_678 (
  .O(mux_o_678),
  .I0(mux_o_673),
  .I1(mux_o_674),
  .S0(dff_q_2)
);
MUX2 mux_inst_679 (
  .O(mux_o_679),
  .I0(mux_o_675),
  .I1(mux_o_676),
  .S0(dff_q_1)
);
MUX2 mux_inst_680 (
  .O(mux_o_680),
  .I0(mux_o_677),
  .I1(mux_o_678),
  .S0(dff_q_1)
);
MUX2 mux_inst_681 (
  .O(dout[21]),
  .I0(mux_o_679),
  .I1(mux_o_680),
  .S0(dff_q_0)
);
MUX2 mux_inst_682 (
  .O(mux_o_682),
  .I0(sp_inst_32_dout[22]),
  .I1(sp_inst_33_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_683 (
  .O(mux_o_683),
  .I0(sp_inst_34_dout[22]),
  .I1(sp_inst_35_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_684 (
  .O(mux_o_684),
  .I0(sp_inst_36_dout[22]),
  .I1(sp_inst_37_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_685 (
  .O(mux_o_685),
  .I0(sp_inst_38_dout[22]),
  .I1(sp_inst_39_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_686 (
  .O(mux_o_686),
  .I0(sp_inst_40_dout[22]),
  .I1(sp_inst_41_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_687 (
  .O(mux_o_687),
  .I0(sp_inst_42_dout[22]),
  .I1(sp_inst_43_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_688 (
  .O(mux_o_688),
  .I0(sp_inst_44_dout[22]),
  .I1(sp_inst_45_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_689 (
  .O(mux_o_689),
  .I0(sp_inst_46_dout[22]),
  .I1(sp_inst_47_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_690 (
  .O(mux_o_690),
  .I0(sp_inst_48_dout[22]),
  .I1(sp_inst_49_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_691 (
  .O(mux_o_691),
  .I0(sp_inst_50_dout[22]),
  .I1(sp_inst_51_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_692 (
  .O(mux_o_692),
  .I0(sp_inst_52_dout[22]),
  .I1(sp_inst_53_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_693 (
  .O(mux_o_693),
  .I0(sp_inst_54_dout[22]),
  .I1(sp_inst_55_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_694 (
  .O(mux_o_694),
  .I0(sp_inst_56_dout[22]),
  .I1(sp_inst_57_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_695 (
  .O(mux_o_695),
  .I0(sp_inst_58_dout[22]),
  .I1(sp_inst_59_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_696 (
  .O(mux_o_696),
  .I0(sp_inst_60_dout[22]),
  .I1(sp_inst_61_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_697 (
  .O(mux_o_697),
  .I0(sp_inst_62_dout[22]),
  .I1(sp_inst_63_dout[22]),
  .S0(dff_q_4)
);
MUX2 mux_inst_698 (
  .O(mux_o_698),
  .I0(mux_o_682),
  .I1(mux_o_683),
  .S0(dff_q_3)
);
MUX2 mux_inst_699 (
  .O(mux_o_699),
  .I0(mux_o_684),
  .I1(mux_o_685),
  .S0(dff_q_3)
);
MUX2 mux_inst_700 (
  .O(mux_o_700),
  .I0(mux_o_686),
  .I1(mux_o_687),
  .S0(dff_q_3)
);
MUX2 mux_inst_701 (
  .O(mux_o_701),
  .I0(mux_o_688),
  .I1(mux_o_689),
  .S0(dff_q_3)
);
MUX2 mux_inst_702 (
  .O(mux_o_702),
  .I0(mux_o_690),
  .I1(mux_o_691),
  .S0(dff_q_3)
);
MUX2 mux_inst_703 (
  .O(mux_o_703),
  .I0(mux_o_692),
  .I1(mux_o_693),
  .S0(dff_q_3)
);
MUX2 mux_inst_704 (
  .O(mux_o_704),
  .I0(mux_o_694),
  .I1(mux_o_695),
  .S0(dff_q_3)
);
MUX2 mux_inst_705 (
  .O(mux_o_705),
  .I0(mux_o_696),
  .I1(mux_o_697),
  .S0(dff_q_3)
);
MUX2 mux_inst_706 (
  .O(mux_o_706),
  .I0(mux_o_698),
  .I1(mux_o_699),
  .S0(dff_q_2)
);
MUX2 mux_inst_707 (
  .O(mux_o_707),
  .I0(mux_o_700),
  .I1(mux_o_701),
  .S0(dff_q_2)
);
MUX2 mux_inst_708 (
  .O(mux_o_708),
  .I0(mux_o_702),
  .I1(mux_o_703),
  .S0(dff_q_2)
);
MUX2 mux_inst_709 (
  .O(mux_o_709),
  .I0(mux_o_704),
  .I1(mux_o_705),
  .S0(dff_q_2)
);
MUX2 mux_inst_710 (
  .O(mux_o_710),
  .I0(mux_o_706),
  .I1(mux_o_707),
  .S0(dff_q_1)
);
MUX2 mux_inst_711 (
  .O(mux_o_711),
  .I0(mux_o_708),
  .I1(mux_o_709),
  .S0(dff_q_1)
);
MUX2 mux_inst_712 (
  .O(dout[22]),
  .I0(mux_o_710),
  .I1(mux_o_711),
  .S0(dff_q_0)
);
MUX2 mux_inst_713 (
  .O(mux_o_713),
  .I0(sp_inst_32_dout[23]),
  .I1(sp_inst_33_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_714 (
  .O(mux_o_714),
  .I0(sp_inst_34_dout[23]),
  .I1(sp_inst_35_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_715 (
  .O(mux_o_715),
  .I0(sp_inst_36_dout[23]),
  .I1(sp_inst_37_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_716 (
  .O(mux_o_716),
  .I0(sp_inst_38_dout[23]),
  .I1(sp_inst_39_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_717 (
  .O(mux_o_717),
  .I0(sp_inst_40_dout[23]),
  .I1(sp_inst_41_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_718 (
  .O(mux_o_718),
  .I0(sp_inst_42_dout[23]),
  .I1(sp_inst_43_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_719 (
  .O(mux_o_719),
  .I0(sp_inst_44_dout[23]),
  .I1(sp_inst_45_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_720 (
  .O(mux_o_720),
  .I0(sp_inst_46_dout[23]),
  .I1(sp_inst_47_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_721 (
  .O(mux_o_721),
  .I0(sp_inst_48_dout[23]),
  .I1(sp_inst_49_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_722 (
  .O(mux_o_722),
  .I0(sp_inst_50_dout[23]),
  .I1(sp_inst_51_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_723 (
  .O(mux_o_723),
  .I0(sp_inst_52_dout[23]),
  .I1(sp_inst_53_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_724 (
  .O(mux_o_724),
  .I0(sp_inst_54_dout[23]),
  .I1(sp_inst_55_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_725 (
  .O(mux_o_725),
  .I0(sp_inst_56_dout[23]),
  .I1(sp_inst_57_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_726 (
  .O(mux_o_726),
  .I0(sp_inst_58_dout[23]),
  .I1(sp_inst_59_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_727 (
  .O(mux_o_727),
  .I0(sp_inst_60_dout[23]),
  .I1(sp_inst_61_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_728 (
  .O(mux_o_728),
  .I0(sp_inst_62_dout[23]),
  .I1(sp_inst_63_dout[23]),
  .S0(dff_q_4)
);
MUX2 mux_inst_729 (
  .O(mux_o_729),
  .I0(mux_o_713),
  .I1(mux_o_714),
  .S0(dff_q_3)
);
MUX2 mux_inst_730 (
  .O(mux_o_730),
  .I0(mux_o_715),
  .I1(mux_o_716),
  .S0(dff_q_3)
);
MUX2 mux_inst_731 (
  .O(mux_o_731),
  .I0(mux_o_717),
  .I1(mux_o_718),
  .S0(dff_q_3)
);
MUX2 mux_inst_732 (
  .O(mux_o_732),
  .I0(mux_o_719),
  .I1(mux_o_720),
  .S0(dff_q_3)
);
MUX2 mux_inst_733 (
  .O(mux_o_733),
  .I0(mux_o_721),
  .I1(mux_o_722),
  .S0(dff_q_3)
);
MUX2 mux_inst_734 (
  .O(mux_o_734),
  .I0(mux_o_723),
  .I1(mux_o_724),
  .S0(dff_q_3)
);
MUX2 mux_inst_735 (
  .O(mux_o_735),
  .I0(mux_o_725),
  .I1(mux_o_726),
  .S0(dff_q_3)
);
MUX2 mux_inst_736 (
  .O(mux_o_736),
  .I0(mux_o_727),
  .I1(mux_o_728),
  .S0(dff_q_3)
);
MUX2 mux_inst_737 (
  .O(mux_o_737),
  .I0(mux_o_729),
  .I1(mux_o_730),
  .S0(dff_q_2)
);
MUX2 mux_inst_738 (
  .O(mux_o_738),
  .I0(mux_o_731),
  .I1(mux_o_732),
  .S0(dff_q_2)
);
MUX2 mux_inst_739 (
  .O(mux_o_739),
  .I0(mux_o_733),
  .I1(mux_o_734),
  .S0(dff_q_2)
);
MUX2 mux_inst_740 (
  .O(mux_o_740),
  .I0(mux_o_735),
  .I1(mux_o_736),
  .S0(dff_q_2)
);
MUX2 mux_inst_741 (
  .O(mux_o_741),
  .I0(mux_o_737),
  .I1(mux_o_738),
  .S0(dff_q_1)
);
MUX2 mux_inst_742 (
  .O(mux_o_742),
  .I0(mux_o_739),
  .I1(mux_o_740),
  .S0(dff_q_1)
);
MUX2 mux_inst_743 (
  .O(dout[23]),
  .I0(mux_o_741),
  .I1(mux_o_742),
  .S0(dff_q_0)
);
MUX2 mux_inst_744 (
  .O(mux_o_744),
  .I0(sp_inst_32_dout[24]),
  .I1(sp_inst_33_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_745 (
  .O(mux_o_745),
  .I0(sp_inst_34_dout[24]),
  .I1(sp_inst_35_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_746 (
  .O(mux_o_746),
  .I0(sp_inst_36_dout[24]),
  .I1(sp_inst_37_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_747 (
  .O(mux_o_747),
  .I0(sp_inst_38_dout[24]),
  .I1(sp_inst_39_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_748 (
  .O(mux_o_748),
  .I0(sp_inst_40_dout[24]),
  .I1(sp_inst_41_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_749 (
  .O(mux_o_749),
  .I0(sp_inst_42_dout[24]),
  .I1(sp_inst_43_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_750 (
  .O(mux_o_750),
  .I0(sp_inst_44_dout[24]),
  .I1(sp_inst_45_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_751 (
  .O(mux_o_751),
  .I0(sp_inst_46_dout[24]),
  .I1(sp_inst_47_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_752 (
  .O(mux_o_752),
  .I0(sp_inst_48_dout[24]),
  .I1(sp_inst_49_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_753 (
  .O(mux_o_753),
  .I0(sp_inst_50_dout[24]),
  .I1(sp_inst_51_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_754 (
  .O(mux_o_754),
  .I0(sp_inst_52_dout[24]),
  .I1(sp_inst_53_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_755 (
  .O(mux_o_755),
  .I0(sp_inst_54_dout[24]),
  .I1(sp_inst_55_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_756 (
  .O(mux_o_756),
  .I0(sp_inst_56_dout[24]),
  .I1(sp_inst_57_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_757 (
  .O(mux_o_757),
  .I0(sp_inst_58_dout[24]),
  .I1(sp_inst_59_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_758 (
  .O(mux_o_758),
  .I0(sp_inst_60_dout[24]),
  .I1(sp_inst_61_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_759 (
  .O(mux_o_759),
  .I0(sp_inst_62_dout[24]),
  .I1(sp_inst_63_dout[24]),
  .S0(dff_q_4)
);
MUX2 mux_inst_760 (
  .O(mux_o_760),
  .I0(mux_o_744),
  .I1(mux_o_745),
  .S0(dff_q_3)
);
MUX2 mux_inst_761 (
  .O(mux_o_761),
  .I0(mux_o_746),
  .I1(mux_o_747),
  .S0(dff_q_3)
);
MUX2 mux_inst_762 (
  .O(mux_o_762),
  .I0(mux_o_748),
  .I1(mux_o_749),
  .S0(dff_q_3)
);
MUX2 mux_inst_763 (
  .O(mux_o_763),
  .I0(mux_o_750),
  .I1(mux_o_751),
  .S0(dff_q_3)
);
MUX2 mux_inst_764 (
  .O(mux_o_764),
  .I0(mux_o_752),
  .I1(mux_o_753),
  .S0(dff_q_3)
);
MUX2 mux_inst_765 (
  .O(mux_o_765),
  .I0(mux_o_754),
  .I1(mux_o_755),
  .S0(dff_q_3)
);
MUX2 mux_inst_766 (
  .O(mux_o_766),
  .I0(mux_o_756),
  .I1(mux_o_757),
  .S0(dff_q_3)
);
MUX2 mux_inst_767 (
  .O(mux_o_767),
  .I0(mux_o_758),
  .I1(mux_o_759),
  .S0(dff_q_3)
);
MUX2 mux_inst_768 (
  .O(mux_o_768),
  .I0(mux_o_760),
  .I1(mux_o_761),
  .S0(dff_q_2)
);
MUX2 mux_inst_769 (
  .O(mux_o_769),
  .I0(mux_o_762),
  .I1(mux_o_763),
  .S0(dff_q_2)
);
MUX2 mux_inst_770 (
  .O(mux_o_770),
  .I0(mux_o_764),
  .I1(mux_o_765),
  .S0(dff_q_2)
);
MUX2 mux_inst_771 (
  .O(mux_o_771),
  .I0(mux_o_766),
  .I1(mux_o_767),
  .S0(dff_q_2)
);
MUX2 mux_inst_772 (
  .O(mux_o_772),
  .I0(mux_o_768),
  .I1(mux_o_769),
  .S0(dff_q_1)
);
MUX2 mux_inst_773 (
  .O(mux_o_773),
  .I0(mux_o_770),
  .I1(mux_o_771),
  .S0(dff_q_1)
);
MUX2 mux_inst_774 (
  .O(dout[24]),
  .I0(mux_o_772),
  .I1(mux_o_773),
  .S0(dff_q_0)
);
MUX2 mux_inst_775 (
  .O(mux_o_775),
  .I0(sp_inst_32_dout[25]),
  .I1(sp_inst_33_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_776 (
  .O(mux_o_776),
  .I0(sp_inst_34_dout[25]),
  .I1(sp_inst_35_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_777 (
  .O(mux_o_777),
  .I0(sp_inst_36_dout[25]),
  .I1(sp_inst_37_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_778 (
  .O(mux_o_778),
  .I0(sp_inst_38_dout[25]),
  .I1(sp_inst_39_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_779 (
  .O(mux_o_779),
  .I0(sp_inst_40_dout[25]),
  .I1(sp_inst_41_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_780 (
  .O(mux_o_780),
  .I0(sp_inst_42_dout[25]),
  .I1(sp_inst_43_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_781 (
  .O(mux_o_781),
  .I0(sp_inst_44_dout[25]),
  .I1(sp_inst_45_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_782 (
  .O(mux_o_782),
  .I0(sp_inst_46_dout[25]),
  .I1(sp_inst_47_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_783 (
  .O(mux_o_783),
  .I0(sp_inst_48_dout[25]),
  .I1(sp_inst_49_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_784 (
  .O(mux_o_784),
  .I0(sp_inst_50_dout[25]),
  .I1(sp_inst_51_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_785 (
  .O(mux_o_785),
  .I0(sp_inst_52_dout[25]),
  .I1(sp_inst_53_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_786 (
  .O(mux_o_786),
  .I0(sp_inst_54_dout[25]),
  .I1(sp_inst_55_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_787 (
  .O(mux_o_787),
  .I0(sp_inst_56_dout[25]),
  .I1(sp_inst_57_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_788 (
  .O(mux_o_788),
  .I0(sp_inst_58_dout[25]),
  .I1(sp_inst_59_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_789 (
  .O(mux_o_789),
  .I0(sp_inst_60_dout[25]),
  .I1(sp_inst_61_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_790 (
  .O(mux_o_790),
  .I0(sp_inst_62_dout[25]),
  .I1(sp_inst_63_dout[25]),
  .S0(dff_q_4)
);
MUX2 mux_inst_791 (
  .O(mux_o_791),
  .I0(mux_o_775),
  .I1(mux_o_776),
  .S0(dff_q_3)
);
MUX2 mux_inst_792 (
  .O(mux_o_792),
  .I0(mux_o_777),
  .I1(mux_o_778),
  .S0(dff_q_3)
);
MUX2 mux_inst_793 (
  .O(mux_o_793),
  .I0(mux_o_779),
  .I1(mux_o_780),
  .S0(dff_q_3)
);
MUX2 mux_inst_794 (
  .O(mux_o_794),
  .I0(mux_o_781),
  .I1(mux_o_782),
  .S0(dff_q_3)
);
MUX2 mux_inst_795 (
  .O(mux_o_795),
  .I0(mux_o_783),
  .I1(mux_o_784),
  .S0(dff_q_3)
);
MUX2 mux_inst_796 (
  .O(mux_o_796),
  .I0(mux_o_785),
  .I1(mux_o_786),
  .S0(dff_q_3)
);
MUX2 mux_inst_797 (
  .O(mux_o_797),
  .I0(mux_o_787),
  .I1(mux_o_788),
  .S0(dff_q_3)
);
MUX2 mux_inst_798 (
  .O(mux_o_798),
  .I0(mux_o_789),
  .I1(mux_o_790),
  .S0(dff_q_3)
);
MUX2 mux_inst_799 (
  .O(mux_o_799),
  .I0(mux_o_791),
  .I1(mux_o_792),
  .S0(dff_q_2)
);
MUX2 mux_inst_800 (
  .O(mux_o_800),
  .I0(mux_o_793),
  .I1(mux_o_794),
  .S0(dff_q_2)
);
MUX2 mux_inst_801 (
  .O(mux_o_801),
  .I0(mux_o_795),
  .I1(mux_o_796),
  .S0(dff_q_2)
);
MUX2 mux_inst_802 (
  .O(mux_o_802),
  .I0(mux_o_797),
  .I1(mux_o_798),
  .S0(dff_q_2)
);
MUX2 mux_inst_803 (
  .O(mux_o_803),
  .I0(mux_o_799),
  .I1(mux_o_800),
  .S0(dff_q_1)
);
MUX2 mux_inst_804 (
  .O(mux_o_804),
  .I0(mux_o_801),
  .I1(mux_o_802),
  .S0(dff_q_1)
);
MUX2 mux_inst_805 (
  .O(dout[25]),
  .I0(mux_o_803),
  .I1(mux_o_804),
  .S0(dff_q_0)
);
MUX2 mux_inst_806 (
  .O(mux_o_806),
  .I0(sp_inst_32_dout[26]),
  .I1(sp_inst_33_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_807 (
  .O(mux_o_807),
  .I0(sp_inst_34_dout[26]),
  .I1(sp_inst_35_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_808 (
  .O(mux_o_808),
  .I0(sp_inst_36_dout[26]),
  .I1(sp_inst_37_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_809 (
  .O(mux_o_809),
  .I0(sp_inst_38_dout[26]),
  .I1(sp_inst_39_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_810 (
  .O(mux_o_810),
  .I0(sp_inst_40_dout[26]),
  .I1(sp_inst_41_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_811 (
  .O(mux_o_811),
  .I0(sp_inst_42_dout[26]),
  .I1(sp_inst_43_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_812 (
  .O(mux_o_812),
  .I0(sp_inst_44_dout[26]),
  .I1(sp_inst_45_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_813 (
  .O(mux_o_813),
  .I0(sp_inst_46_dout[26]),
  .I1(sp_inst_47_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_814 (
  .O(mux_o_814),
  .I0(sp_inst_48_dout[26]),
  .I1(sp_inst_49_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_815 (
  .O(mux_o_815),
  .I0(sp_inst_50_dout[26]),
  .I1(sp_inst_51_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_816 (
  .O(mux_o_816),
  .I0(sp_inst_52_dout[26]),
  .I1(sp_inst_53_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_817 (
  .O(mux_o_817),
  .I0(sp_inst_54_dout[26]),
  .I1(sp_inst_55_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_818 (
  .O(mux_o_818),
  .I0(sp_inst_56_dout[26]),
  .I1(sp_inst_57_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_819 (
  .O(mux_o_819),
  .I0(sp_inst_58_dout[26]),
  .I1(sp_inst_59_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_820 (
  .O(mux_o_820),
  .I0(sp_inst_60_dout[26]),
  .I1(sp_inst_61_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_821 (
  .O(mux_o_821),
  .I0(sp_inst_62_dout[26]),
  .I1(sp_inst_63_dout[26]),
  .S0(dff_q_4)
);
MUX2 mux_inst_822 (
  .O(mux_o_822),
  .I0(mux_o_806),
  .I1(mux_o_807),
  .S0(dff_q_3)
);
MUX2 mux_inst_823 (
  .O(mux_o_823),
  .I0(mux_o_808),
  .I1(mux_o_809),
  .S0(dff_q_3)
);
MUX2 mux_inst_824 (
  .O(mux_o_824),
  .I0(mux_o_810),
  .I1(mux_o_811),
  .S0(dff_q_3)
);
MUX2 mux_inst_825 (
  .O(mux_o_825),
  .I0(mux_o_812),
  .I1(mux_o_813),
  .S0(dff_q_3)
);
MUX2 mux_inst_826 (
  .O(mux_o_826),
  .I0(mux_o_814),
  .I1(mux_o_815),
  .S0(dff_q_3)
);
MUX2 mux_inst_827 (
  .O(mux_o_827),
  .I0(mux_o_816),
  .I1(mux_o_817),
  .S0(dff_q_3)
);
MUX2 mux_inst_828 (
  .O(mux_o_828),
  .I0(mux_o_818),
  .I1(mux_o_819),
  .S0(dff_q_3)
);
MUX2 mux_inst_829 (
  .O(mux_o_829),
  .I0(mux_o_820),
  .I1(mux_o_821),
  .S0(dff_q_3)
);
MUX2 mux_inst_830 (
  .O(mux_o_830),
  .I0(mux_o_822),
  .I1(mux_o_823),
  .S0(dff_q_2)
);
MUX2 mux_inst_831 (
  .O(mux_o_831),
  .I0(mux_o_824),
  .I1(mux_o_825),
  .S0(dff_q_2)
);
MUX2 mux_inst_832 (
  .O(mux_o_832),
  .I0(mux_o_826),
  .I1(mux_o_827),
  .S0(dff_q_2)
);
MUX2 mux_inst_833 (
  .O(mux_o_833),
  .I0(mux_o_828),
  .I1(mux_o_829),
  .S0(dff_q_2)
);
MUX2 mux_inst_834 (
  .O(mux_o_834),
  .I0(mux_o_830),
  .I1(mux_o_831),
  .S0(dff_q_1)
);
MUX2 mux_inst_835 (
  .O(mux_o_835),
  .I0(mux_o_832),
  .I1(mux_o_833),
  .S0(dff_q_1)
);
MUX2 mux_inst_836 (
  .O(dout[26]),
  .I0(mux_o_834),
  .I1(mux_o_835),
  .S0(dff_q_0)
);
MUX2 mux_inst_837 (
  .O(mux_o_837),
  .I0(sp_inst_32_dout[27]),
  .I1(sp_inst_33_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_838 (
  .O(mux_o_838),
  .I0(sp_inst_34_dout[27]),
  .I1(sp_inst_35_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_839 (
  .O(mux_o_839),
  .I0(sp_inst_36_dout[27]),
  .I1(sp_inst_37_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_840 (
  .O(mux_o_840),
  .I0(sp_inst_38_dout[27]),
  .I1(sp_inst_39_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_841 (
  .O(mux_o_841),
  .I0(sp_inst_40_dout[27]),
  .I1(sp_inst_41_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_842 (
  .O(mux_o_842),
  .I0(sp_inst_42_dout[27]),
  .I1(sp_inst_43_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_843 (
  .O(mux_o_843),
  .I0(sp_inst_44_dout[27]),
  .I1(sp_inst_45_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_844 (
  .O(mux_o_844),
  .I0(sp_inst_46_dout[27]),
  .I1(sp_inst_47_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_845 (
  .O(mux_o_845),
  .I0(sp_inst_48_dout[27]),
  .I1(sp_inst_49_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_846 (
  .O(mux_o_846),
  .I0(sp_inst_50_dout[27]),
  .I1(sp_inst_51_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_847 (
  .O(mux_o_847),
  .I0(sp_inst_52_dout[27]),
  .I1(sp_inst_53_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_848 (
  .O(mux_o_848),
  .I0(sp_inst_54_dout[27]),
  .I1(sp_inst_55_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_849 (
  .O(mux_o_849),
  .I0(sp_inst_56_dout[27]),
  .I1(sp_inst_57_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_850 (
  .O(mux_o_850),
  .I0(sp_inst_58_dout[27]),
  .I1(sp_inst_59_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_851 (
  .O(mux_o_851),
  .I0(sp_inst_60_dout[27]),
  .I1(sp_inst_61_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_852 (
  .O(mux_o_852),
  .I0(sp_inst_62_dout[27]),
  .I1(sp_inst_63_dout[27]),
  .S0(dff_q_4)
);
MUX2 mux_inst_853 (
  .O(mux_o_853),
  .I0(mux_o_837),
  .I1(mux_o_838),
  .S0(dff_q_3)
);
MUX2 mux_inst_854 (
  .O(mux_o_854),
  .I0(mux_o_839),
  .I1(mux_o_840),
  .S0(dff_q_3)
);
MUX2 mux_inst_855 (
  .O(mux_o_855),
  .I0(mux_o_841),
  .I1(mux_o_842),
  .S0(dff_q_3)
);
MUX2 mux_inst_856 (
  .O(mux_o_856),
  .I0(mux_o_843),
  .I1(mux_o_844),
  .S0(dff_q_3)
);
MUX2 mux_inst_857 (
  .O(mux_o_857),
  .I0(mux_o_845),
  .I1(mux_o_846),
  .S0(dff_q_3)
);
MUX2 mux_inst_858 (
  .O(mux_o_858),
  .I0(mux_o_847),
  .I1(mux_o_848),
  .S0(dff_q_3)
);
MUX2 mux_inst_859 (
  .O(mux_o_859),
  .I0(mux_o_849),
  .I1(mux_o_850),
  .S0(dff_q_3)
);
MUX2 mux_inst_860 (
  .O(mux_o_860),
  .I0(mux_o_851),
  .I1(mux_o_852),
  .S0(dff_q_3)
);
MUX2 mux_inst_861 (
  .O(mux_o_861),
  .I0(mux_o_853),
  .I1(mux_o_854),
  .S0(dff_q_2)
);
MUX2 mux_inst_862 (
  .O(mux_o_862),
  .I0(mux_o_855),
  .I1(mux_o_856),
  .S0(dff_q_2)
);
MUX2 mux_inst_863 (
  .O(mux_o_863),
  .I0(mux_o_857),
  .I1(mux_o_858),
  .S0(dff_q_2)
);
MUX2 mux_inst_864 (
  .O(mux_o_864),
  .I0(mux_o_859),
  .I1(mux_o_860),
  .S0(dff_q_2)
);
MUX2 mux_inst_865 (
  .O(mux_o_865),
  .I0(mux_o_861),
  .I1(mux_o_862),
  .S0(dff_q_1)
);
MUX2 mux_inst_866 (
  .O(mux_o_866),
  .I0(mux_o_863),
  .I1(mux_o_864),
  .S0(dff_q_1)
);
MUX2 mux_inst_867 (
  .O(dout[27]),
  .I0(mux_o_865),
  .I1(mux_o_866),
  .S0(dff_q_0)
);
MUX2 mux_inst_868 (
  .O(mux_o_868),
  .I0(sp_inst_32_dout[28]),
  .I1(sp_inst_33_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_869 (
  .O(mux_o_869),
  .I0(sp_inst_34_dout[28]),
  .I1(sp_inst_35_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_870 (
  .O(mux_o_870),
  .I0(sp_inst_36_dout[28]),
  .I1(sp_inst_37_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_871 (
  .O(mux_o_871),
  .I0(sp_inst_38_dout[28]),
  .I1(sp_inst_39_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_872 (
  .O(mux_o_872),
  .I0(sp_inst_40_dout[28]),
  .I1(sp_inst_41_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_873 (
  .O(mux_o_873),
  .I0(sp_inst_42_dout[28]),
  .I1(sp_inst_43_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_874 (
  .O(mux_o_874),
  .I0(sp_inst_44_dout[28]),
  .I1(sp_inst_45_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_875 (
  .O(mux_o_875),
  .I0(sp_inst_46_dout[28]),
  .I1(sp_inst_47_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_876 (
  .O(mux_o_876),
  .I0(sp_inst_48_dout[28]),
  .I1(sp_inst_49_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_877 (
  .O(mux_o_877),
  .I0(sp_inst_50_dout[28]),
  .I1(sp_inst_51_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_878 (
  .O(mux_o_878),
  .I0(sp_inst_52_dout[28]),
  .I1(sp_inst_53_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_879 (
  .O(mux_o_879),
  .I0(sp_inst_54_dout[28]),
  .I1(sp_inst_55_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_880 (
  .O(mux_o_880),
  .I0(sp_inst_56_dout[28]),
  .I1(sp_inst_57_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_881 (
  .O(mux_o_881),
  .I0(sp_inst_58_dout[28]),
  .I1(sp_inst_59_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_882 (
  .O(mux_o_882),
  .I0(sp_inst_60_dout[28]),
  .I1(sp_inst_61_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_883 (
  .O(mux_o_883),
  .I0(sp_inst_62_dout[28]),
  .I1(sp_inst_63_dout[28]),
  .S0(dff_q_4)
);
MUX2 mux_inst_884 (
  .O(mux_o_884),
  .I0(mux_o_868),
  .I1(mux_o_869),
  .S0(dff_q_3)
);
MUX2 mux_inst_885 (
  .O(mux_o_885),
  .I0(mux_o_870),
  .I1(mux_o_871),
  .S0(dff_q_3)
);
MUX2 mux_inst_886 (
  .O(mux_o_886),
  .I0(mux_o_872),
  .I1(mux_o_873),
  .S0(dff_q_3)
);
MUX2 mux_inst_887 (
  .O(mux_o_887),
  .I0(mux_o_874),
  .I1(mux_o_875),
  .S0(dff_q_3)
);
MUX2 mux_inst_888 (
  .O(mux_o_888),
  .I0(mux_o_876),
  .I1(mux_o_877),
  .S0(dff_q_3)
);
MUX2 mux_inst_889 (
  .O(mux_o_889),
  .I0(mux_o_878),
  .I1(mux_o_879),
  .S0(dff_q_3)
);
MUX2 mux_inst_890 (
  .O(mux_o_890),
  .I0(mux_o_880),
  .I1(mux_o_881),
  .S0(dff_q_3)
);
MUX2 mux_inst_891 (
  .O(mux_o_891),
  .I0(mux_o_882),
  .I1(mux_o_883),
  .S0(dff_q_3)
);
MUX2 mux_inst_892 (
  .O(mux_o_892),
  .I0(mux_o_884),
  .I1(mux_o_885),
  .S0(dff_q_2)
);
MUX2 mux_inst_893 (
  .O(mux_o_893),
  .I0(mux_o_886),
  .I1(mux_o_887),
  .S0(dff_q_2)
);
MUX2 mux_inst_894 (
  .O(mux_o_894),
  .I0(mux_o_888),
  .I1(mux_o_889),
  .S0(dff_q_2)
);
MUX2 mux_inst_895 (
  .O(mux_o_895),
  .I0(mux_o_890),
  .I1(mux_o_891),
  .S0(dff_q_2)
);
MUX2 mux_inst_896 (
  .O(mux_o_896),
  .I0(mux_o_892),
  .I1(mux_o_893),
  .S0(dff_q_1)
);
MUX2 mux_inst_897 (
  .O(mux_o_897),
  .I0(mux_o_894),
  .I1(mux_o_895),
  .S0(dff_q_1)
);
MUX2 mux_inst_898 (
  .O(dout[28]),
  .I0(mux_o_896),
  .I1(mux_o_897),
  .S0(dff_q_0)
);
MUX2 mux_inst_899 (
  .O(mux_o_899),
  .I0(sp_inst_32_dout[29]),
  .I1(sp_inst_33_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_900 (
  .O(mux_o_900),
  .I0(sp_inst_34_dout[29]),
  .I1(sp_inst_35_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_901 (
  .O(mux_o_901),
  .I0(sp_inst_36_dout[29]),
  .I1(sp_inst_37_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_902 (
  .O(mux_o_902),
  .I0(sp_inst_38_dout[29]),
  .I1(sp_inst_39_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_903 (
  .O(mux_o_903),
  .I0(sp_inst_40_dout[29]),
  .I1(sp_inst_41_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_904 (
  .O(mux_o_904),
  .I0(sp_inst_42_dout[29]),
  .I1(sp_inst_43_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_905 (
  .O(mux_o_905),
  .I0(sp_inst_44_dout[29]),
  .I1(sp_inst_45_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_906 (
  .O(mux_o_906),
  .I0(sp_inst_46_dout[29]),
  .I1(sp_inst_47_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_907 (
  .O(mux_o_907),
  .I0(sp_inst_48_dout[29]),
  .I1(sp_inst_49_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_908 (
  .O(mux_o_908),
  .I0(sp_inst_50_dout[29]),
  .I1(sp_inst_51_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_909 (
  .O(mux_o_909),
  .I0(sp_inst_52_dout[29]),
  .I1(sp_inst_53_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_910 (
  .O(mux_o_910),
  .I0(sp_inst_54_dout[29]),
  .I1(sp_inst_55_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_911 (
  .O(mux_o_911),
  .I0(sp_inst_56_dout[29]),
  .I1(sp_inst_57_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_912 (
  .O(mux_o_912),
  .I0(sp_inst_58_dout[29]),
  .I1(sp_inst_59_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_913 (
  .O(mux_o_913),
  .I0(sp_inst_60_dout[29]),
  .I1(sp_inst_61_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_914 (
  .O(mux_o_914),
  .I0(sp_inst_62_dout[29]),
  .I1(sp_inst_63_dout[29]),
  .S0(dff_q_4)
);
MUX2 mux_inst_915 (
  .O(mux_o_915),
  .I0(mux_o_899),
  .I1(mux_o_900),
  .S0(dff_q_3)
);
MUX2 mux_inst_916 (
  .O(mux_o_916),
  .I0(mux_o_901),
  .I1(mux_o_902),
  .S0(dff_q_3)
);
MUX2 mux_inst_917 (
  .O(mux_o_917),
  .I0(mux_o_903),
  .I1(mux_o_904),
  .S0(dff_q_3)
);
MUX2 mux_inst_918 (
  .O(mux_o_918),
  .I0(mux_o_905),
  .I1(mux_o_906),
  .S0(dff_q_3)
);
MUX2 mux_inst_919 (
  .O(mux_o_919),
  .I0(mux_o_907),
  .I1(mux_o_908),
  .S0(dff_q_3)
);
MUX2 mux_inst_920 (
  .O(mux_o_920),
  .I0(mux_o_909),
  .I1(mux_o_910),
  .S0(dff_q_3)
);
MUX2 mux_inst_921 (
  .O(mux_o_921),
  .I0(mux_o_911),
  .I1(mux_o_912),
  .S0(dff_q_3)
);
MUX2 mux_inst_922 (
  .O(mux_o_922),
  .I0(mux_o_913),
  .I1(mux_o_914),
  .S0(dff_q_3)
);
MUX2 mux_inst_923 (
  .O(mux_o_923),
  .I0(mux_o_915),
  .I1(mux_o_916),
  .S0(dff_q_2)
);
MUX2 mux_inst_924 (
  .O(mux_o_924),
  .I0(mux_o_917),
  .I1(mux_o_918),
  .S0(dff_q_2)
);
MUX2 mux_inst_925 (
  .O(mux_o_925),
  .I0(mux_o_919),
  .I1(mux_o_920),
  .S0(dff_q_2)
);
MUX2 mux_inst_926 (
  .O(mux_o_926),
  .I0(mux_o_921),
  .I1(mux_o_922),
  .S0(dff_q_2)
);
MUX2 mux_inst_927 (
  .O(mux_o_927),
  .I0(mux_o_923),
  .I1(mux_o_924),
  .S0(dff_q_1)
);
MUX2 mux_inst_928 (
  .O(mux_o_928),
  .I0(mux_o_925),
  .I1(mux_o_926),
  .S0(dff_q_1)
);
MUX2 mux_inst_929 (
  .O(dout[29]),
  .I0(mux_o_927),
  .I1(mux_o_928),
  .S0(dff_q_0)
);
MUX2 mux_inst_930 (
  .O(mux_o_930),
  .I0(sp_inst_32_dout[30]),
  .I1(sp_inst_33_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_931 (
  .O(mux_o_931),
  .I0(sp_inst_34_dout[30]),
  .I1(sp_inst_35_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_932 (
  .O(mux_o_932),
  .I0(sp_inst_36_dout[30]),
  .I1(sp_inst_37_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_933 (
  .O(mux_o_933),
  .I0(sp_inst_38_dout[30]),
  .I1(sp_inst_39_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_934 (
  .O(mux_o_934),
  .I0(sp_inst_40_dout[30]),
  .I1(sp_inst_41_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_935 (
  .O(mux_o_935),
  .I0(sp_inst_42_dout[30]),
  .I1(sp_inst_43_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_936 (
  .O(mux_o_936),
  .I0(sp_inst_44_dout[30]),
  .I1(sp_inst_45_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_937 (
  .O(mux_o_937),
  .I0(sp_inst_46_dout[30]),
  .I1(sp_inst_47_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_938 (
  .O(mux_o_938),
  .I0(sp_inst_48_dout[30]),
  .I1(sp_inst_49_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_939 (
  .O(mux_o_939),
  .I0(sp_inst_50_dout[30]),
  .I1(sp_inst_51_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_940 (
  .O(mux_o_940),
  .I0(sp_inst_52_dout[30]),
  .I1(sp_inst_53_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_941 (
  .O(mux_o_941),
  .I0(sp_inst_54_dout[30]),
  .I1(sp_inst_55_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_942 (
  .O(mux_o_942),
  .I0(sp_inst_56_dout[30]),
  .I1(sp_inst_57_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_943 (
  .O(mux_o_943),
  .I0(sp_inst_58_dout[30]),
  .I1(sp_inst_59_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_944 (
  .O(mux_o_944),
  .I0(sp_inst_60_dout[30]),
  .I1(sp_inst_61_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_945 (
  .O(mux_o_945),
  .I0(sp_inst_62_dout[30]),
  .I1(sp_inst_63_dout[30]),
  .S0(dff_q_4)
);
MUX2 mux_inst_946 (
  .O(mux_o_946),
  .I0(mux_o_930),
  .I1(mux_o_931),
  .S0(dff_q_3)
);
MUX2 mux_inst_947 (
  .O(mux_o_947),
  .I0(mux_o_932),
  .I1(mux_o_933),
  .S0(dff_q_3)
);
MUX2 mux_inst_948 (
  .O(mux_o_948),
  .I0(mux_o_934),
  .I1(mux_o_935),
  .S0(dff_q_3)
);
MUX2 mux_inst_949 (
  .O(mux_o_949),
  .I0(mux_o_936),
  .I1(mux_o_937),
  .S0(dff_q_3)
);
MUX2 mux_inst_950 (
  .O(mux_o_950),
  .I0(mux_o_938),
  .I1(mux_o_939),
  .S0(dff_q_3)
);
MUX2 mux_inst_951 (
  .O(mux_o_951),
  .I0(mux_o_940),
  .I1(mux_o_941),
  .S0(dff_q_3)
);
MUX2 mux_inst_952 (
  .O(mux_o_952),
  .I0(mux_o_942),
  .I1(mux_o_943),
  .S0(dff_q_3)
);
MUX2 mux_inst_953 (
  .O(mux_o_953),
  .I0(mux_o_944),
  .I1(mux_o_945),
  .S0(dff_q_3)
);
MUX2 mux_inst_954 (
  .O(mux_o_954),
  .I0(mux_o_946),
  .I1(mux_o_947),
  .S0(dff_q_2)
);
MUX2 mux_inst_955 (
  .O(mux_o_955),
  .I0(mux_o_948),
  .I1(mux_o_949),
  .S0(dff_q_2)
);
MUX2 mux_inst_956 (
  .O(mux_o_956),
  .I0(mux_o_950),
  .I1(mux_o_951),
  .S0(dff_q_2)
);
MUX2 mux_inst_957 (
  .O(mux_o_957),
  .I0(mux_o_952),
  .I1(mux_o_953),
  .S0(dff_q_2)
);
MUX2 mux_inst_958 (
  .O(mux_o_958),
  .I0(mux_o_954),
  .I1(mux_o_955),
  .S0(dff_q_1)
);
MUX2 mux_inst_959 (
  .O(mux_o_959),
  .I0(mux_o_956),
  .I1(mux_o_957),
  .S0(dff_q_1)
);
MUX2 mux_inst_960 (
  .O(dout[30]),
  .I0(mux_o_958),
  .I1(mux_o_959),
  .S0(dff_q_0)
);
MUX2 mux_inst_961 (
  .O(mux_o_961),
  .I0(sp_inst_32_dout[31]),
  .I1(sp_inst_33_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_962 (
  .O(mux_o_962),
  .I0(sp_inst_34_dout[31]),
  .I1(sp_inst_35_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_963 (
  .O(mux_o_963),
  .I0(sp_inst_36_dout[31]),
  .I1(sp_inst_37_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_964 (
  .O(mux_o_964),
  .I0(sp_inst_38_dout[31]),
  .I1(sp_inst_39_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_965 (
  .O(mux_o_965),
  .I0(sp_inst_40_dout[31]),
  .I1(sp_inst_41_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_966 (
  .O(mux_o_966),
  .I0(sp_inst_42_dout[31]),
  .I1(sp_inst_43_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_967 (
  .O(mux_o_967),
  .I0(sp_inst_44_dout[31]),
  .I1(sp_inst_45_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_968 (
  .O(mux_o_968),
  .I0(sp_inst_46_dout[31]),
  .I1(sp_inst_47_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_969 (
  .O(mux_o_969),
  .I0(sp_inst_48_dout[31]),
  .I1(sp_inst_49_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_970 (
  .O(mux_o_970),
  .I0(sp_inst_50_dout[31]),
  .I1(sp_inst_51_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_971 (
  .O(mux_o_971),
  .I0(sp_inst_52_dout[31]),
  .I1(sp_inst_53_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_972 (
  .O(mux_o_972),
  .I0(sp_inst_54_dout[31]),
  .I1(sp_inst_55_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_973 (
  .O(mux_o_973),
  .I0(sp_inst_56_dout[31]),
  .I1(sp_inst_57_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_974 (
  .O(mux_o_974),
  .I0(sp_inst_58_dout[31]),
  .I1(sp_inst_59_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_975 (
  .O(mux_o_975),
  .I0(sp_inst_60_dout[31]),
  .I1(sp_inst_61_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_976 (
  .O(mux_o_976),
  .I0(sp_inst_62_dout[31]),
  .I1(sp_inst_63_dout[31]),
  .S0(dff_q_4)
);
MUX2 mux_inst_977 (
  .O(mux_o_977),
  .I0(mux_o_961),
  .I1(mux_o_962),
  .S0(dff_q_3)
);
MUX2 mux_inst_978 (
  .O(mux_o_978),
  .I0(mux_o_963),
  .I1(mux_o_964),
  .S0(dff_q_3)
);
MUX2 mux_inst_979 (
  .O(mux_o_979),
  .I0(mux_o_965),
  .I1(mux_o_966),
  .S0(dff_q_3)
);
MUX2 mux_inst_980 (
  .O(mux_o_980),
  .I0(mux_o_967),
  .I1(mux_o_968),
  .S0(dff_q_3)
);
MUX2 mux_inst_981 (
  .O(mux_o_981),
  .I0(mux_o_969),
  .I1(mux_o_970),
  .S0(dff_q_3)
);
MUX2 mux_inst_982 (
  .O(mux_o_982),
  .I0(mux_o_971),
  .I1(mux_o_972),
  .S0(dff_q_3)
);
MUX2 mux_inst_983 (
  .O(mux_o_983),
  .I0(mux_o_973),
  .I1(mux_o_974),
  .S0(dff_q_3)
);
MUX2 mux_inst_984 (
  .O(mux_o_984),
  .I0(mux_o_975),
  .I1(mux_o_976),
  .S0(dff_q_3)
);
MUX2 mux_inst_985 (
  .O(mux_o_985),
  .I0(mux_o_977),
  .I1(mux_o_978),
  .S0(dff_q_2)
);
MUX2 mux_inst_986 (
  .O(mux_o_986),
  .I0(mux_o_979),
  .I1(mux_o_980),
  .S0(dff_q_2)
);
MUX2 mux_inst_987 (
  .O(mux_o_987),
  .I0(mux_o_981),
  .I1(mux_o_982),
  .S0(dff_q_2)
);
MUX2 mux_inst_988 (
  .O(mux_o_988),
  .I0(mux_o_983),
  .I1(mux_o_984),
  .S0(dff_q_2)
);
MUX2 mux_inst_989 (
  .O(mux_o_989),
  .I0(mux_o_985),
  .I1(mux_o_986),
  .S0(dff_q_1)
);
MUX2 mux_inst_990 (
  .O(mux_o_990),
  .I0(mux_o_987),
  .I1(mux_o_988),
  .S0(dff_q_1)
);
MUX2 mux_inst_991 (
  .O(dout[31]),
  .I0(mux_o_989),
  .I1(mux_o_990),
  .S0(dff_q_0)
);
endmodule //blk_mem_gen_0
